module rol(
  input         clock,
  input         reset,
  input  [31:0] io_num,
  input  [31:0] io_cnt,
  input         io_valid,
  output        io_ready,
  output [31:0] io_out_rol
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[rol.scala 14:24]
  wire [1:0] _GEN_0 = reset ? 2'h3 : state; // @[rol.scala 15:26 16:15 14:24]
  reg [31:0] temp; // @[rol.scala 18:19]
  wire [1:0] _state_T = io_valid ? 2'h0 : state; // @[rol.scala 23:25]
  wire [31:0] _temp_T = io_cnt; // @[rol.scala 26:47]
  wire [62:0] _GEN_10 = {{31{io_num[31]}},io_num}; // @[rol.scala 26:29]
  wire [62:0] _temp_T_2 = $signed(_GEN_10) << _temp_T[4:0]; // @[rol.scala 26:29]
  wire [31:0] _temp_T_7 = 32'sh20 - $signed(io_cnt); // @[rol.scala 30:77]
  wire [31:0] _temp_T_10 = io_num >> _temp_T_7[4:0]; // @[rol.scala 30:92]
  wire [31:0] _temp_T_12 = $signed(temp) | $signed(_temp_T_10); // @[rol.scala 30:26]
  wire [2:0] _GEN_1 = 2'h2 == state ? 3'h7 : {{1'd0}, _GEN_0}; // @[rol.scala 21:19 34:19]
  wire [31:0] _GEN_2 = 2'h1 == state ? $signed(_temp_T_12) : $signed(temp); // @[rol.scala 21:19 30:18 18:19]
  wire [2:0] _GEN_3 = 2'h1 == state ? 3'h2 : _GEN_1; // @[rol.scala 21:19 31:19]
  wire [62:0] _GEN_4 = 2'h0 == state ? $signed(_temp_T_2) : $signed({{31{_GEN_2[31]}},_GEN_2}); // @[rol.scala 21:19 26:18]
  wire [2:0] _GEN_5 = 2'h0 == state ? 3'h1 : _GEN_3; // @[rol.scala 21:19 27:19]
  wire [2:0] _GEN_6 = 2'h3 == state ? {{1'd0}, _state_T} : _GEN_5; // @[rol.scala 21:19 23:19]
  wire [62:0] _GEN_7 = 2'h3 == state ? $signed({{31{temp[31]}},temp}) : $signed(_GEN_4); // @[rol.scala 18:19 21:19]
  wire [2:0] _GEN_8 = reset ? 3'h3 : _GEN_6; // @[rol.scala 14:{24,24}]
  assign io_ready = state == 2'h2; // @[rol.scala 38:23]
  assign io_out_rol = temp; // @[rol.scala 19:16]
  always @(posedge clock) begin
    state <= _GEN_8[1:0]; // @[rol.scala 14:{24,24}]
    temp <= _GEN_7[31:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  temp = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module fill(
  input         clock,
  input         reset,
  input  [31:0] io_value,
  input  [31:0] io_arr_0,
  input  [31:0] io_arr_1,
  input  [31:0] io_arr_2,
  input  [31:0] io_arr_3,
  input  [31:0] io_arr_4,
  input  [31:0] io_arr_5,
  input  [31:0] io_arr_6,
  input  [31:0] io_arr_7,
  input  [31:0] io_arr_8,
  input  [31:0] io_arr_9,
  input  [31:0] io_arr_10,
  input  [31:0] io_arr_11,
  input  [31:0] io_arr_12,
  input  [31:0] io_arr_13,
  input  [31:0] io_arr_14,
  input  [31:0] io_arr_15,
  input  [31:0] io_arr_16,
  input  [31:0] io_arr_17,
  input  [31:0] io_arr_18,
  input  [31:0] io_arr_19,
  input  [31:0] io_arr_20,
  input  [31:0] io_arr_21,
  input  [31:0] io_arr_22,
  input  [31:0] io_arr_23,
  input  [31:0] io_arr_24,
  input  [31:0] io_arr_25,
  input  [31:0] io_arr_26,
  input  [31:0] io_arr_27,
  input  [31:0] io_arr_28,
  input  [31:0] io_arr_29,
  input  [31:0] io_arr_30,
  input  [31:0] io_arr_31,
  input  [31:0] io_arr_32,
  input  [31:0] io_arr_33,
  input  [31:0] io_arr_34,
  input  [31:0] io_arr_35,
  input  [31:0] io_arr_36,
  input  [31:0] io_arr_37,
  input  [31:0] io_arr_38,
  input  [31:0] io_arr_39,
  input  [31:0] io_arr_40,
  input  [31:0] io_arr_41,
  input  [31:0] io_arr_42,
  input  [31:0] io_arr_43,
  input  [31:0] io_arr_44,
  input  [31:0] io_arr_45,
  input  [31:0] io_arr_46,
  input  [31:0] io_arr_47,
  input  [31:0] io_arr_48,
  input  [31:0] io_arr_49,
  input  [31:0] io_arr_50,
  input  [31:0] io_arr_51,
  input  [31:0] io_arr_52,
  input  [31:0] io_arr_53,
  input  [31:0] io_arr_54,
  input  [31:0] io_arr_55,
  input  [31:0] io_arr_56,
  input  [31:0] io_arr_57,
  input  [31:0] io_arr_58,
  input  [31:0] io_arr_59,
  input  [31:0] io_arr_60,
  input  [31:0] io_arr_61,
  input  [31:0] io_arr_62,
  input  [31:0] io_arr_63,
  input  [31:0] io_arr_64,
  input  [31:0] io_arr_65,
  input  [31:0] io_arr_66,
  input  [31:0] io_arr_67,
  input  [31:0] io_arr_68,
  input  [31:0] io_arr_69,
  input  [31:0] io_arr_70,
  input  [31:0] io_arr_71,
  input  [31:0] io_arr_72,
  input  [31:0] io_arr_73,
  input  [31:0] io_arr_74,
  input  [31:0] io_arr_75,
  input  [31:0] io_arr_76,
  input  [31:0] io_arr_77,
  input  [31:0] io_arr_78,
  input  [31:0] io_arr_79,
  input  [31:0] io_off,
  input         io_valid,
  output [31:0] io_arr_out_0,
  output [31:0] io_arr_out_1,
  output [31:0] io_arr_out_2,
  output [31:0] io_arr_out_3,
  output [31:0] io_arr_out_4,
  output [31:0] io_arr_out_5,
  output [31:0] io_arr_out_6,
  output [31:0] io_arr_out_7,
  output [31:0] io_arr_out_8,
  output [31:0] io_arr_out_9,
  output [31:0] io_arr_out_10,
  output [31:0] io_arr_out_11,
  output [31:0] io_arr_out_12,
  output [31:0] io_arr_out_13,
  output [31:0] io_arr_out_14,
  output [31:0] io_arr_out_15,
  output [31:0] io_arr_out_16,
  output [31:0] io_arr_out_17,
  output [31:0] io_arr_out_18,
  output [31:0] io_arr_out_19,
  output [31:0] io_arr_out_20,
  output [31:0] io_arr_out_21,
  output [31:0] io_arr_out_22,
  output [31:0] io_arr_out_23,
  output [31:0] io_arr_out_24,
  output [31:0] io_arr_out_25,
  output [31:0] io_arr_out_26,
  output [31:0] io_arr_out_27,
  output [31:0] io_arr_out_28,
  output [31:0] io_arr_out_29,
  output [31:0] io_arr_out_30,
  output [31:0] io_arr_out_31,
  output [31:0] io_arr_out_32,
  output [31:0] io_arr_out_33,
  output [31:0] io_arr_out_34,
  output [31:0] io_arr_out_35,
  output [31:0] io_arr_out_36,
  output [31:0] io_arr_out_37,
  output [31:0] io_arr_out_38,
  output [31:0] io_arr_out_39,
  output [31:0] io_arr_out_40,
  output [31:0] io_arr_out_41,
  output [31:0] io_arr_out_42,
  output [31:0] io_arr_out_43,
  output [31:0] io_arr_out_44,
  output [31:0] io_arr_out_45,
  output [31:0] io_arr_out_46,
  output [31:0] io_arr_out_47,
  output [31:0] io_arr_out_48,
  output [31:0] io_arr_out_49,
  output [31:0] io_arr_out_50,
  output [31:0] io_arr_out_51,
  output [31:0] io_arr_out_52,
  output [31:0] io_arr_out_53,
  output [31:0] io_arr_out_54,
  output [31:0] io_arr_out_55,
  output [31:0] io_arr_out_56,
  output [31:0] io_arr_out_57,
  output [31:0] io_arr_out_58,
  output [31:0] io_arr_out_59,
  output [31:0] io_arr_out_60,
  output [31:0] io_arr_out_61,
  output [31:0] io_arr_out_62,
  output [31:0] io_arr_out_63,
  output [31:0] io_arr_out_64,
  output [31:0] io_arr_out_65,
  output [31:0] io_arr_out_66,
  output [31:0] io_arr_out_67,
  output [31:0] io_arr_out_68,
  output [31:0] io_arr_out_69,
  output [31:0] io_arr_out_70,
  output [31:0] io_arr_out_71,
  output [31:0] io_arr_out_72,
  output [31:0] io_arr_out_73,
  output [31:0] io_arr_out_74,
  output [31:0] io_arr_out_75,
  output [31:0] io_arr_out_76,
  output [31:0] io_arr_out_77,
  output [31:0] io_arr_out_78,
  output [31:0] io_arr_out_79,
  output        io_ready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[fill.scala 15:24]
  wire [2:0] _GEN_0 = reset ? 3'h7 : state; // @[fill.scala 16:26 17:15 15:24]
  reg [31:0] arr_0; // @[fill.scala 19:18]
  reg [31:0] arr_1; // @[fill.scala 19:18]
  reg [31:0] arr_2; // @[fill.scala 19:18]
  reg [31:0] arr_3; // @[fill.scala 19:18]
  reg [31:0] arr_4; // @[fill.scala 19:18]
  reg [31:0] arr_5; // @[fill.scala 19:18]
  reg [31:0] arr_6; // @[fill.scala 19:18]
  reg [31:0] arr_7; // @[fill.scala 19:18]
  reg [31:0] arr_8; // @[fill.scala 19:18]
  reg [31:0] arr_9; // @[fill.scala 19:18]
  reg [31:0] arr_10; // @[fill.scala 19:18]
  reg [31:0] arr_11; // @[fill.scala 19:18]
  reg [31:0] arr_12; // @[fill.scala 19:18]
  reg [31:0] arr_13; // @[fill.scala 19:18]
  reg [31:0] arr_14; // @[fill.scala 19:18]
  reg [31:0] arr_15; // @[fill.scala 19:18]
  reg [31:0] arr_16; // @[fill.scala 19:18]
  reg [31:0] arr_17; // @[fill.scala 19:18]
  reg [31:0] arr_18; // @[fill.scala 19:18]
  reg [31:0] arr_19; // @[fill.scala 19:18]
  reg [31:0] arr_20; // @[fill.scala 19:18]
  reg [31:0] arr_21; // @[fill.scala 19:18]
  reg [31:0] arr_22; // @[fill.scala 19:18]
  reg [31:0] arr_23; // @[fill.scala 19:18]
  reg [31:0] arr_24; // @[fill.scala 19:18]
  reg [31:0] arr_25; // @[fill.scala 19:18]
  reg [31:0] arr_26; // @[fill.scala 19:18]
  reg [31:0] arr_27; // @[fill.scala 19:18]
  reg [31:0] arr_28; // @[fill.scala 19:18]
  reg [31:0] arr_29; // @[fill.scala 19:18]
  reg [31:0] arr_30; // @[fill.scala 19:18]
  reg [31:0] arr_31; // @[fill.scala 19:18]
  reg [31:0] arr_32; // @[fill.scala 19:18]
  reg [31:0] arr_33; // @[fill.scala 19:18]
  reg [31:0] arr_34; // @[fill.scala 19:18]
  reg [31:0] arr_35; // @[fill.scala 19:18]
  reg [31:0] arr_36; // @[fill.scala 19:18]
  reg [31:0] arr_37; // @[fill.scala 19:18]
  reg [31:0] arr_38; // @[fill.scala 19:18]
  reg [31:0] arr_39; // @[fill.scala 19:18]
  reg [31:0] arr_40; // @[fill.scala 19:18]
  reg [31:0] arr_41; // @[fill.scala 19:18]
  reg [31:0] arr_42; // @[fill.scala 19:18]
  reg [31:0] arr_43; // @[fill.scala 19:18]
  reg [31:0] arr_44; // @[fill.scala 19:18]
  reg [31:0] arr_45; // @[fill.scala 19:18]
  reg [31:0] arr_46; // @[fill.scala 19:18]
  reg [31:0] arr_47; // @[fill.scala 19:18]
  reg [31:0] arr_48; // @[fill.scala 19:18]
  reg [31:0] arr_49; // @[fill.scala 19:18]
  reg [31:0] arr_50; // @[fill.scala 19:18]
  reg [31:0] arr_51; // @[fill.scala 19:18]
  reg [31:0] arr_52; // @[fill.scala 19:18]
  reg [31:0] arr_53; // @[fill.scala 19:18]
  reg [31:0] arr_54; // @[fill.scala 19:18]
  reg [31:0] arr_55; // @[fill.scala 19:18]
  reg [31:0] arr_56; // @[fill.scala 19:18]
  reg [31:0] arr_57; // @[fill.scala 19:18]
  reg [31:0] arr_58; // @[fill.scala 19:18]
  reg [31:0] arr_59; // @[fill.scala 19:18]
  reg [31:0] arr_60; // @[fill.scala 19:18]
  reg [31:0] arr_61; // @[fill.scala 19:18]
  reg [31:0] arr_62; // @[fill.scala 19:18]
  reg [31:0] arr_63; // @[fill.scala 19:18]
  reg [31:0] arr_64; // @[fill.scala 19:18]
  reg [31:0] arr_65; // @[fill.scala 19:18]
  reg [31:0] arr_66; // @[fill.scala 19:18]
  reg [31:0] arr_67; // @[fill.scala 19:18]
  reg [31:0] arr_68; // @[fill.scala 19:18]
  reg [31:0] arr_69; // @[fill.scala 19:18]
  reg [31:0] arr_70; // @[fill.scala 19:18]
  reg [31:0] arr_71; // @[fill.scala 19:18]
  reg [31:0] arr_72; // @[fill.scala 19:18]
  reg [31:0] arr_73; // @[fill.scala 19:18]
  reg [31:0] arr_74; // @[fill.scala 19:18]
  reg [31:0] arr_75; // @[fill.scala 19:18]
  reg [31:0] arr_76; // @[fill.scala 19:18]
  reg [31:0] arr_77; // @[fill.scala 19:18]
  reg [31:0] arr_78; // @[fill.scala 19:18]
  reg [31:0] arr_79; // @[fill.scala 19:18]
  reg  REG; // @[fill.scala 20:17]
  wire [31:0] _GEN_1 = REG ? $signed(io_arr_0) : $signed(arr_0); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_2 = REG ? $signed(io_arr_1) : $signed(arr_1); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_3 = REG ? $signed(io_arr_2) : $signed(arr_2); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_4 = REG ? $signed(io_arr_3) : $signed(arr_3); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_5 = REG ? $signed(io_arr_4) : $signed(arr_4); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_6 = REG ? $signed(io_arr_5) : $signed(arr_5); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_7 = REG ? $signed(io_arr_6) : $signed(arr_6); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_8 = REG ? $signed(io_arr_7) : $signed(arr_7); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_9 = REG ? $signed(io_arr_8) : $signed(arr_8); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_10 = REG ? $signed(io_arr_9) : $signed(arr_9); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_11 = REG ? $signed(io_arr_10) : $signed(arr_10); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_12 = REG ? $signed(io_arr_11) : $signed(arr_11); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_13 = REG ? $signed(io_arr_12) : $signed(arr_12); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_14 = REG ? $signed(io_arr_13) : $signed(arr_13); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_15 = REG ? $signed(io_arr_14) : $signed(arr_14); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_16 = REG ? $signed(io_arr_15) : $signed(arr_15); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_17 = REG ? $signed(io_arr_16) : $signed(arr_16); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_18 = REG ? $signed(io_arr_17) : $signed(arr_17); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_19 = REG ? $signed(io_arr_18) : $signed(arr_18); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_20 = REG ? $signed(io_arr_19) : $signed(arr_19); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_21 = REG ? $signed(io_arr_20) : $signed(arr_20); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_22 = REG ? $signed(io_arr_21) : $signed(arr_21); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_23 = REG ? $signed(io_arr_22) : $signed(arr_22); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_24 = REG ? $signed(io_arr_23) : $signed(arr_23); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_25 = REG ? $signed(io_arr_24) : $signed(arr_24); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_26 = REG ? $signed(io_arr_25) : $signed(arr_25); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_27 = REG ? $signed(io_arr_26) : $signed(arr_26); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_28 = REG ? $signed(io_arr_27) : $signed(arr_27); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_29 = REG ? $signed(io_arr_28) : $signed(arr_28); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_30 = REG ? $signed(io_arr_29) : $signed(arr_29); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_31 = REG ? $signed(io_arr_30) : $signed(arr_30); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_32 = REG ? $signed(io_arr_31) : $signed(arr_31); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_33 = REG ? $signed(io_arr_32) : $signed(arr_32); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_34 = REG ? $signed(io_arr_33) : $signed(arr_33); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_35 = REG ? $signed(io_arr_34) : $signed(arr_34); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_36 = REG ? $signed(io_arr_35) : $signed(arr_35); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_37 = REG ? $signed(io_arr_36) : $signed(arr_36); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_38 = REG ? $signed(io_arr_37) : $signed(arr_37); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_39 = REG ? $signed(io_arr_38) : $signed(arr_38); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_40 = REG ? $signed(io_arr_39) : $signed(arr_39); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_41 = REG ? $signed(io_arr_40) : $signed(arr_40); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_42 = REG ? $signed(io_arr_41) : $signed(arr_41); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_43 = REG ? $signed(io_arr_42) : $signed(arr_42); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_44 = REG ? $signed(io_arr_43) : $signed(arr_43); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_45 = REG ? $signed(io_arr_44) : $signed(arr_44); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_46 = REG ? $signed(io_arr_45) : $signed(arr_45); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_47 = REG ? $signed(io_arr_46) : $signed(arr_46); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_48 = REG ? $signed(io_arr_47) : $signed(arr_47); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_49 = REG ? $signed(io_arr_48) : $signed(arr_48); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_50 = REG ? $signed(io_arr_49) : $signed(arr_49); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_51 = REG ? $signed(io_arr_50) : $signed(arr_50); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_52 = REG ? $signed(io_arr_51) : $signed(arr_51); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_53 = REG ? $signed(io_arr_52) : $signed(arr_52); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_54 = REG ? $signed(io_arr_53) : $signed(arr_53); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_55 = REG ? $signed(io_arr_54) : $signed(arr_54); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_56 = REG ? $signed(io_arr_55) : $signed(arr_55); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_57 = REG ? $signed(io_arr_56) : $signed(arr_56); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_58 = REG ? $signed(io_arr_57) : $signed(arr_57); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_59 = REG ? $signed(io_arr_58) : $signed(arr_58); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_60 = REG ? $signed(io_arr_59) : $signed(arr_59); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_61 = REG ? $signed(io_arr_60) : $signed(arr_60); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_62 = REG ? $signed(io_arr_61) : $signed(arr_61); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_63 = REG ? $signed(io_arr_62) : $signed(arr_62); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_64 = REG ? $signed(io_arr_63) : $signed(arr_63); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_65 = REG ? $signed(io_arr_64) : $signed(arr_64); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_66 = REG ? $signed(io_arr_65) : $signed(arr_65); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_67 = REG ? $signed(io_arr_66) : $signed(arr_66); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_68 = REG ? $signed(io_arr_67) : $signed(arr_67); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_69 = REG ? $signed(io_arr_68) : $signed(arr_68); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_70 = REG ? $signed(io_arr_69) : $signed(arr_69); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_71 = REG ? $signed(io_arr_70) : $signed(arr_70); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_72 = REG ? $signed(io_arr_71) : $signed(arr_71); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_73 = REG ? $signed(io_arr_72) : $signed(arr_72); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_74 = REG ? $signed(io_arr_73) : $signed(arr_73); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_75 = REG ? $signed(io_arr_74) : $signed(arr_74); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_76 = REG ? $signed(io_arr_75) : $signed(arr_75); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_77 = REG ? $signed(io_arr_76) : $signed(arr_76); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_78 = REG ? $signed(io_arr_77) : $signed(arr_77); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_79 = REG ? $signed(io_arr_78) : $signed(arr_78); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _GEN_80 = REG ? $signed(io_arr_79) : $signed(arr_79); // @[fill.scala 20:29 21:13 19:18]
  wire [31:0] _T_4 = io_off; // @[fill.scala 30:32]
  wire [31:0] _arr_T = io_value; // @[fill.scala 30:55]
  wire [31:0] _arr_T_4 = {{24'd0}, _arr_T[31:24]}; // @[fill.scala 30:96]
  wire [31:0] _arr_T_6 = $signed(_arr_T_4) & 32'shff; // @[fill.scala 30:99]
  wire [31:0] _T_10 = $signed(io_off) + 32'sh1; // @[fill.scala 34:45]
  wire [31:0] _arr_T_11 = {{16'd0}, _arr_T[31:16]}; // @[fill.scala 34:109]
  wire [31:0] _arr_T_13 = $signed(_arr_T_11) & 32'shff; // @[fill.scala 34:112]
  wire [31:0] _T_16 = $signed(io_off) + 32'sh2; // @[fill.scala 38:45]
  wire [31:0] _arr_T_18 = {{8'd0}, _arr_T[31:8]}; // @[fill.scala 38:108]
  wire [31:0] _arr_T_20 = $signed(_arr_T_18) & 32'shff; // @[fill.scala 38:111]
  wire [31:0] _GEN_241 = 7'h0 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_1); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_242 = 7'h1 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_2); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_243 = 7'h2 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_3); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_244 = 7'h3 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_4); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_245 = 7'h4 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_5); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_246 = 7'h5 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_6); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_247 = 7'h6 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_7); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_248 = 7'h7 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_8); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_249 = 7'h8 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_9); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_250 = 7'h9 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_10); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_251 = 7'ha == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_11); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_252 = 7'hb == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_12); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_253 = 7'hc == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_13); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_254 = 7'hd == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_14); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_255 = 7'he == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_15); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_256 = 7'hf == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_16); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_257 = 7'h10 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_17); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_258 = 7'h11 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_18); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_259 = 7'h12 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_19); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_260 = 7'h13 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_20); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_261 = 7'h14 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_21); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_262 = 7'h15 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_22); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_263 = 7'h16 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_23); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_264 = 7'h17 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_24); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_265 = 7'h18 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_25); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_266 = 7'h19 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_26); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_267 = 7'h1a == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_27); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_268 = 7'h1b == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_28); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_269 = 7'h1c == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_29); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_270 = 7'h1d == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_30); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_271 = 7'h1e == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_31); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_272 = 7'h1f == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_32); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_273 = 7'h20 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_33); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_274 = 7'h21 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_34); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_275 = 7'h22 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_35); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_276 = 7'h23 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_36); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_277 = 7'h24 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_37); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_278 = 7'h25 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_38); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_279 = 7'h26 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_39); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_280 = 7'h27 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_40); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_281 = 7'h28 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_41); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_282 = 7'h29 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_42); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_283 = 7'h2a == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_43); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_284 = 7'h2b == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_44); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_285 = 7'h2c == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_45); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_286 = 7'h2d == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_46); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_287 = 7'h2e == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_47); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_288 = 7'h2f == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_48); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_289 = 7'h30 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_49); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_290 = 7'h31 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_50); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_291 = 7'h32 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_51); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_292 = 7'h33 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_52); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_293 = 7'h34 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_53); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_294 = 7'h35 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_54); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_295 = 7'h36 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_55); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_296 = 7'h37 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_56); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_297 = 7'h38 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_57); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_298 = 7'h39 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_58); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_299 = 7'h3a == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_59); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_300 = 7'h3b == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_60); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_301 = 7'h3c == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_61); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_302 = 7'h3d == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_62); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_303 = 7'h3e == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_63); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_304 = 7'h3f == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_64); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_305 = 7'h40 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_65); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_306 = 7'h41 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_66); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_307 = 7'h42 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_67); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_308 = 7'h43 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_68); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_309 = 7'h44 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_69); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_310 = 7'h45 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_70); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_311 = 7'h46 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_71); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_312 = 7'h47 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_72); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_313 = 7'h48 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_73); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_314 = 7'h49 == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_74); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_315 = 7'h4a == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_75); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_316 = 7'h4b == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_76); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_317 = 7'h4c == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_77); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_318 = 7'h4d == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_78); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_319 = 7'h4e == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_79); // @[fill.scala 38:{49,49}]
  wire [31:0] _GEN_320 = 7'h4f == _T_16[6:0] ? $signed(_arr_T_20) : $signed(_GEN_80); // @[fill.scala 38:{49,49}]
  wire [31:0] _T_22 = $signed(io_off) + 32'sh3; // @[fill.scala 42:45]
  wire [31:0] _arr_T_22 = $signed(io_value) & 32'shff; // @[fill.scala 42:61]
  wire [31:0] _GEN_321 = 7'h0 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_1); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_322 = 7'h1 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_2); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_323 = 7'h2 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_3); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_324 = 7'h3 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_4); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_325 = 7'h4 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_5); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_326 = 7'h5 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_6); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_327 = 7'h6 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_7); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_328 = 7'h7 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_8); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_329 = 7'h8 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_9); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_330 = 7'h9 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_10); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_331 = 7'ha == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_11); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_332 = 7'hb == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_12); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_333 = 7'hc == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_13); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_334 = 7'hd == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_14); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_335 = 7'he == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_15); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_336 = 7'hf == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_16); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_337 = 7'h10 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_17); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_338 = 7'h11 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_18); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_339 = 7'h12 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_19); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_340 = 7'h13 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_20); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_341 = 7'h14 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_21); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_342 = 7'h15 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_22); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_343 = 7'h16 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_23); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_344 = 7'h17 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_24); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_345 = 7'h18 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_25); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_346 = 7'h19 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_26); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_347 = 7'h1a == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_27); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_348 = 7'h1b == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_28); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_349 = 7'h1c == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_29); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_350 = 7'h1d == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_30); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_351 = 7'h1e == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_31); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_352 = 7'h1f == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_32); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_353 = 7'h20 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_33); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_354 = 7'h21 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_34); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_355 = 7'h22 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_35); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_356 = 7'h23 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_36); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_357 = 7'h24 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_37); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_358 = 7'h25 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_38); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_359 = 7'h26 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_39); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_360 = 7'h27 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_40); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_361 = 7'h28 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_41); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_362 = 7'h29 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_42); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_363 = 7'h2a == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_43); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_364 = 7'h2b == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_44); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_365 = 7'h2c == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_45); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_366 = 7'h2d == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_46); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_367 = 7'h2e == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_47); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_368 = 7'h2f == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_48); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_369 = 7'h30 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_49); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_370 = 7'h31 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_50); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_371 = 7'h32 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_51); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_372 = 7'h33 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_52); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_373 = 7'h34 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_53); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_374 = 7'h35 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_54); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_375 = 7'h36 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_55); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_376 = 7'h37 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_56); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_377 = 7'h38 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_57); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_378 = 7'h39 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_58); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_379 = 7'h3a == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_59); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_380 = 7'h3b == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_60); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_381 = 7'h3c == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_61); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_382 = 7'h3d == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_62); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_383 = 7'h3e == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_63); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_384 = 7'h3f == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_64); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_385 = 7'h40 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_65); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_386 = 7'h41 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_66); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_387 = 7'h42 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_67); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_388 = 7'h43 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_68); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_389 = 7'h44 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_69); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_390 = 7'h45 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_70); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_391 = 7'h46 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_71); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_392 = 7'h47 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_72); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_393 = 7'h48 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_73); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_394 = 7'h49 == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_74); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_395 = 7'h4a == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_75); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_396 = 7'h4b == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_76); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_397 = 7'h4c == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_77); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_398 = 7'h4d == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_78); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_399 = 7'h4e == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_79); // @[fill.scala 42:{49,49}]
  wire [31:0] _GEN_400 = 7'h4f == _T_22[6:0] ? $signed(_arr_T_22) : $signed(_GEN_80); // @[fill.scala 42:{49,49}]
  wire [2:0] _GEN_401 = 3'h4 == state ? 3'h7 : _GEN_0; // @[fill.scala 25:19 46:19]
  wire [31:0] _GEN_402 = 3'h3 == state ? $signed(_GEN_321) : $signed(_GEN_1); // @[fill.scala 25:19]
  wire [31:0] _GEN_403 = 3'h3 == state ? $signed(_GEN_322) : $signed(_GEN_2); // @[fill.scala 25:19]
  wire [31:0] _GEN_404 = 3'h3 == state ? $signed(_GEN_323) : $signed(_GEN_3); // @[fill.scala 25:19]
  wire [31:0] _GEN_405 = 3'h3 == state ? $signed(_GEN_324) : $signed(_GEN_4); // @[fill.scala 25:19]
  wire [31:0] _GEN_406 = 3'h3 == state ? $signed(_GEN_325) : $signed(_GEN_5); // @[fill.scala 25:19]
  wire [31:0] _GEN_407 = 3'h3 == state ? $signed(_GEN_326) : $signed(_GEN_6); // @[fill.scala 25:19]
  wire [31:0] _GEN_408 = 3'h3 == state ? $signed(_GEN_327) : $signed(_GEN_7); // @[fill.scala 25:19]
  wire [31:0] _GEN_409 = 3'h3 == state ? $signed(_GEN_328) : $signed(_GEN_8); // @[fill.scala 25:19]
  wire [31:0] _GEN_410 = 3'h3 == state ? $signed(_GEN_329) : $signed(_GEN_9); // @[fill.scala 25:19]
  wire [31:0] _GEN_411 = 3'h3 == state ? $signed(_GEN_330) : $signed(_GEN_10); // @[fill.scala 25:19]
  wire [31:0] _GEN_412 = 3'h3 == state ? $signed(_GEN_331) : $signed(_GEN_11); // @[fill.scala 25:19]
  wire [31:0] _GEN_413 = 3'h3 == state ? $signed(_GEN_332) : $signed(_GEN_12); // @[fill.scala 25:19]
  wire [31:0] _GEN_414 = 3'h3 == state ? $signed(_GEN_333) : $signed(_GEN_13); // @[fill.scala 25:19]
  wire [31:0] _GEN_415 = 3'h3 == state ? $signed(_GEN_334) : $signed(_GEN_14); // @[fill.scala 25:19]
  wire [31:0] _GEN_416 = 3'h3 == state ? $signed(_GEN_335) : $signed(_GEN_15); // @[fill.scala 25:19]
  wire [31:0] _GEN_417 = 3'h3 == state ? $signed(_GEN_336) : $signed(_GEN_16); // @[fill.scala 25:19]
  wire [31:0] _GEN_418 = 3'h3 == state ? $signed(_GEN_337) : $signed(_GEN_17); // @[fill.scala 25:19]
  wire [31:0] _GEN_419 = 3'h3 == state ? $signed(_GEN_338) : $signed(_GEN_18); // @[fill.scala 25:19]
  wire [31:0] _GEN_420 = 3'h3 == state ? $signed(_GEN_339) : $signed(_GEN_19); // @[fill.scala 25:19]
  wire [31:0] _GEN_421 = 3'h3 == state ? $signed(_GEN_340) : $signed(_GEN_20); // @[fill.scala 25:19]
  wire [31:0] _GEN_422 = 3'h3 == state ? $signed(_GEN_341) : $signed(_GEN_21); // @[fill.scala 25:19]
  wire [31:0] _GEN_423 = 3'h3 == state ? $signed(_GEN_342) : $signed(_GEN_22); // @[fill.scala 25:19]
  wire [31:0] _GEN_424 = 3'h3 == state ? $signed(_GEN_343) : $signed(_GEN_23); // @[fill.scala 25:19]
  wire [31:0] _GEN_425 = 3'h3 == state ? $signed(_GEN_344) : $signed(_GEN_24); // @[fill.scala 25:19]
  wire [31:0] _GEN_426 = 3'h3 == state ? $signed(_GEN_345) : $signed(_GEN_25); // @[fill.scala 25:19]
  wire [31:0] _GEN_427 = 3'h3 == state ? $signed(_GEN_346) : $signed(_GEN_26); // @[fill.scala 25:19]
  wire [31:0] _GEN_428 = 3'h3 == state ? $signed(_GEN_347) : $signed(_GEN_27); // @[fill.scala 25:19]
  wire [31:0] _GEN_429 = 3'h3 == state ? $signed(_GEN_348) : $signed(_GEN_28); // @[fill.scala 25:19]
  wire [31:0] _GEN_430 = 3'h3 == state ? $signed(_GEN_349) : $signed(_GEN_29); // @[fill.scala 25:19]
  wire [31:0] _GEN_431 = 3'h3 == state ? $signed(_GEN_350) : $signed(_GEN_30); // @[fill.scala 25:19]
  wire [31:0] _GEN_432 = 3'h3 == state ? $signed(_GEN_351) : $signed(_GEN_31); // @[fill.scala 25:19]
  wire [31:0] _GEN_433 = 3'h3 == state ? $signed(_GEN_352) : $signed(_GEN_32); // @[fill.scala 25:19]
  wire [31:0] _GEN_434 = 3'h3 == state ? $signed(_GEN_353) : $signed(_GEN_33); // @[fill.scala 25:19]
  wire [31:0] _GEN_435 = 3'h3 == state ? $signed(_GEN_354) : $signed(_GEN_34); // @[fill.scala 25:19]
  wire [31:0] _GEN_436 = 3'h3 == state ? $signed(_GEN_355) : $signed(_GEN_35); // @[fill.scala 25:19]
  wire [31:0] _GEN_437 = 3'h3 == state ? $signed(_GEN_356) : $signed(_GEN_36); // @[fill.scala 25:19]
  wire [31:0] _GEN_438 = 3'h3 == state ? $signed(_GEN_357) : $signed(_GEN_37); // @[fill.scala 25:19]
  wire [31:0] _GEN_439 = 3'h3 == state ? $signed(_GEN_358) : $signed(_GEN_38); // @[fill.scala 25:19]
  wire [31:0] _GEN_440 = 3'h3 == state ? $signed(_GEN_359) : $signed(_GEN_39); // @[fill.scala 25:19]
  wire [31:0] _GEN_441 = 3'h3 == state ? $signed(_GEN_360) : $signed(_GEN_40); // @[fill.scala 25:19]
  wire [31:0] _GEN_442 = 3'h3 == state ? $signed(_GEN_361) : $signed(_GEN_41); // @[fill.scala 25:19]
  wire [31:0] _GEN_443 = 3'h3 == state ? $signed(_GEN_362) : $signed(_GEN_42); // @[fill.scala 25:19]
  wire [31:0] _GEN_444 = 3'h3 == state ? $signed(_GEN_363) : $signed(_GEN_43); // @[fill.scala 25:19]
  wire [31:0] _GEN_445 = 3'h3 == state ? $signed(_GEN_364) : $signed(_GEN_44); // @[fill.scala 25:19]
  wire [31:0] _GEN_446 = 3'h3 == state ? $signed(_GEN_365) : $signed(_GEN_45); // @[fill.scala 25:19]
  wire [31:0] _GEN_447 = 3'h3 == state ? $signed(_GEN_366) : $signed(_GEN_46); // @[fill.scala 25:19]
  wire [31:0] _GEN_448 = 3'h3 == state ? $signed(_GEN_367) : $signed(_GEN_47); // @[fill.scala 25:19]
  wire [31:0] _GEN_449 = 3'h3 == state ? $signed(_GEN_368) : $signed(_GEN_48); // @[fill.scala 25:19]
  wire [31:0] _GEN_450 = 3'h3 == state ? $signed(_GEN_369) : $signed(_GEN_49); // @[fill.scala 25:19]
  wire [31:0] _GEN_451 = 3'h3 == state ? $signed(_GEN_370) : $signed(_GEN_50); // @[fill.scala 25:19]
  wire [31:0] _GEN_452 = 3'h3 == state ? $signed(_GEN_371) : $signed(_GEN_51); // @[fill.scala 25:19]
  wire [31:0] _GEN_453 = 3'h3 == state ? $signed(_GEN_372) : $signed(_GEN_52); // @[fill.scala 25:19]
  wire [31:0] _GEN_454 = 3'h3 == state ? $signed(_GEN_373) : $signed(_GEN_53); // @[fill.scala 25:19]
  wire [31:0] _GEN_455 = 3'h3 == state ? $signed(_GEN_374) : $signed(_GEN_54); // @[fill.scala 25:19]
  wire [31:0] _GEN_456 = 3'h3 == state ? $signed(_GEN_375) : $signed(_GEN_55); // @[fill.scala 25:19]
  wire [31:0] _GEN_457 = 3'h3 == state ? $signed(_GEN_376) : $signed(_GEN_56); // @[fill.scala 25:19]
  wire [31:0] _GEN_458 = 3'h3 == state ? $signed(_GEN_377) : $signed(_GEN_57); // @[fill.scala 25:19]
  wire [31:0] _GEN_459 = 3'h3 == state ? $signed(_GEN_378) : $signed(_GEN_58); // @[fill.scala 25:19]
  wire [31:0] _GEN_460 = 3'h3 == state ? $signed(_GEN_379) : $signed(_GEN_59); // @[fill.scala 25:19]
  wire [31:0] _GEN_461 = 3'h3 == state ? $signed(_GEN_380) : $signed(_GEN_60); // @[fill.scala 25:19]
  wire [31:0] _GEN_462 = 3'h3 == state ? $signed(_GEN_381) : $signed(_GEN_61); // @[fill.scala 25:19]
  wire [31:0] _GEN_463 = 3'h3 == state ? $signed(_GEN_382) : $signed(_GEN_62); // @[fill.scala 25:19]
  wire [31:0] _GEN_464 = 3'h3 == state ? $signed(_GEN_383) : $signed(_GEN_63); // @[fill.scala 25:19]
  wire [31:0] _GEN_465 = 3'h3 == state ? $signed(_GEN_384) : $signed(_GEN_64); // @[fill.scala 25:19]
  wire [31:0] _GEN_466 = 3'h3 == state ? $signed(_GEN_385) : $signed(_GEN_65); // @[fill.scala 25:19]
  wire [31:0] _GEN_467 = 3'h3 == state ? $signed(_GEN_386) : $signed(_GEN_66); // @[fill.scala 25:19]
  wire [31:0] _GEN_468 = 3'h3 == state ? $signed(_GEN_387) : $signed(_GEN_67); // @[fill.scala 25:19]
  wire [31:0] _GEN_469 = 3'h3 == state ? $signed(_GEN_388) : $signed(_GEN_68); // @[fill.scala 25:19]
  wire [31:0] _GEN_470 = 3'h3 == state ? $signed(_GEN_389) : $signed(_GEN_69); // @[fill.scala 25:19]
  wire [31:0] _GEN_471 = 3'h3 == state ? $signed(_GEN_390) : $signed(_GEN_70); // @[fill.scala 25:19]
  wire [31:0] _GEN_472 = 3'h3 == state ? $signed(_GEN_391) : $signed(_GEN_71); // @[fill.scala 25:19]
  wire [31:0] _GEN_473 = 3'h3 == state ? $signed(_GEN_392) : $signed(_GEN_72); // @[fill.scala 25:19]
  wire [31:0] _GEN_474 = 3'h3 == state ? $signed(_GEN_393) : $signed(_GEN_73); // @[fill.scala 25:19]
  wire [31:0] _GEN_475 = 3'h3 == state ? $signed(_GEN_394) : $signed(_GEN_74); // @[fill.scala 25:19]
  wire [31:0] _GEN_476 = 3'h3 == state ? $signed(_GEN_395) : $signed(_GEN_75); // @[fill.scala 25:19]
  wire [31:0] _GEN_477 = 3'h3 == state ? $signed(_GEN_396) : $signed(_GEN_76); // @[fill.scala 25:19]
  wire [31:0] _GEN_478 = 3'h3 == state ? $signed(_GEN_397) : $signed(_GEN_77); // @[fill.scala 25:19]
  wire [31:0] _GEN_479 = 3'h3 == state ? $signed(_GEN_398) : $signed(_GEN_78); // @[fill.scala 25:19]
  wire [31:0] _GEN_480 = 3'h3 == state ? $signed(_GEN_399) : $signed(_GEN_79); // @[fill.scala 25:19]
  wire [31:0] _GEN_481 = 3'h3 == state ? $signed(_GEN_400) : $signed(_GEN_80); // @[fill.scala 25:19]
  wire [2:0] _GEN_482 = 3'h3 == state ? 3'h4 : _GEN_401; // @[fill.scala 25:19 43:19]
  wire [2:0] _GEN_563 = 3'h2 == state ? 3'h3 : _GEN_482; // @[fill.scala 25:19 39:19]
  assign io_arr_out_0 = arr_0; // @[fill.scala 23:16]
  assign io_arr_out_1 = arr_1; // @[fill.scala 23:16]
  assign io_arr_out_2 = arr_2; // @[fill.scala 23:16]
  assign io_arr_out_3 = arr_3; // @[fill.scala 23:16]
  assign io_arr_out_4 = arr_4; // @[fill.scala 23:16]
  assign io_arr_out_5 = arr_5; // @[fill.scala 23:16]
  assign io_arr_out_6 = arr_6; // @[fill.scala 23:16]
  assign io_arr_out_7 = arr_7; // @[fill.scala 23:16]
  assign io_arr_out_8 = arr_8; // @[fill.scala 23:16]
  assign io_arr_out_9 = arr_9; // @[fill.scala 23:16]
  assign io_arr_out_10 = arr_10; // @[fill.scala 23:16]
  assign io_arr_out_11 = arr_11; // @[fill.scala 23:16]
  assign io_arr_out_12 = arr_12; // @[fill.scala 23:16]
  assign io_arr_out_13 = arr_13; // @[fill.scala 23:16]
  assign io_arr_out_14 = arr_14; // @[fill.scala 23:16]
  assign io_arr_out_15 = arr_15; // @[fill.scala 23:16]
  assign io_arr_out_16 = arr_16; // @[fill.scala 23:16]
  assign io_arr_out_17 = arr_17; // @[fill.scala 23:16]
  assign io_arr_out_18 = arr_18; // @[fill.scala 23:16]
  assign io_arr_out_19 = arr_19; // @[fill.scala 23:16]
  assign io_arr_out_20 = arr_20; // @[fill.scala 23:16]
  assign io_arr_out_21 = arr_21; // @[fill.scala 23:16]
  assign io_arr_out_22 = arr_22; // @[fill.scala 23:16]
  assign io_arr_out_23 = arr_23; // @[fill.scala 23:16]
  assign io_arr_out_24 = arr_24; // @[fill.scala 23:16]
  assign io_arr_out_25 = arr_25; // @[fill.scala 23:16]
  assign io_arr_out_26 = arr_26; // @[fill.scala 23:16]
  assign io_arr_out_27 = arr_27; // @[fill.scala 23:16]
  assign io_arr_out_28 = arr_28; // @[fill.scala 23:16]
  assign io_arr_out_29 = arr_29; // @[fill.scala 23:16]
  assign io_arr_out_30 = arr_30; // @[fill.scala 23:16]
  assign io_arr_out_31 = arr_31; // @[fill.scala 23:16]
  assign io_arr_out_32 = arr_32; // @[fill.scala 23:16]
  assign io_arr_out_33 = arr_33; // @[fill.scala 23:16]
  assign io_arr_out_34 = arr_34; // @[fill.scala 23:16]
  assign io_arr_out_35 = arr_35; // @[fill.scala 23:16]
  assign io_arr_out_36 = arr_36; // @[fill.scala 23:16]
  assign io_arr_out_37 = arr_37; // @[fill.scala 23:16]
  assign io_arr_out_38 = arr_38; // @[fill.scala 23:16]
  assign io_arr_out_39 = arr_39; // @[fill.scala 23:16]
  assign io_arr_out_40 = arr_40; // @[fill.scala 23:16]
  assign io_arr_out_41 = arr_41; // @[fill.scala 23:16]
  assign io_arr_out_42 = arr_42; // @[fill.scala 23:16]
  assign io_arr_out_43 = arr_43; // @[fill.scala 23:16]
  assign io_arr_out_44 = arr_44; // @[fill.scala 23:16]
  assign io_arr_out_45 = arr_45; // @[fill.scala 23:16]
  assign io_arr_out_46 = arr_46; // @[fill.scala 23:16]
  assign io_arr_out_47 = arr_47; // @[fill.scala 23:16]
  assign io_arr_out_48 = arr_48; // @[fill.scala 23:16]
  assign io_arr_out_49 = arr_49; // @[fill.scala 23:16]
  assign io_arr_out_50 = arr_50; // @[fill.scala 23:16]
  assign io_arr_out_51 = arr_51; // @[fill.scala 23:16]
  assign io_arr_out_52 = arr_52; // @[fill.scala 23:16]
  assign io_arr_out_53 = arr_53; // @[fill.scala 23:16]
  assign io_arr_out_54 = arr_54; // @[fill.scala 23:16]
  assign io_arr_out_55 = arr_55; // @[fill.scala 23:16]
  assign io_arr_out_56 = arr_56; // @[fill.scala 23:16]
  assign io_arr_out_57 = arr_57; // @[fill.scala 23:16]
  assign io_arr_out_58 = arr_58; // @[fill.scala 23:16]
  assign io_arr_out_59 = arr_59; // @[fill.scala 23:16]
  assign io_arr_out_60 = arr_60; // @[fill.scala 23:16]
  assign io_arr_out_61 = arr_61; // @[fill.scala 23:16]
  assign io_arr_out_62 = arr_62; // @[fill.scala 23:16]
  assign io_arr_out_63 = arr_63; // @[fill.scala 23:16]
  assign io_arr_out_64 = arr_64; // @[fill.scala 23:16]
  assign io_arr_out_65 = arr_65; // @[fill.scala 23:16]
  assign io_arr_out_66 = arr_66; // @[fill.scala 23:16]
  assign io_arr_out_67 = arr_67; // @[fill.scala 23:16]
  assign io_arr_out_68 = arr_68; // @[fill.scala 23:16]
  assign io_arr_out_69 = arr_69; // @[fill.scala 23:16]
  assign io_arr_out_70 = arr_70; // @[fill.scala 23:16]
  assign io_arr_out_71 = arr_71; // @[fill.scala 23:16]
  assign io_arr_out_72 = arr_72; // @[fill.scala 23:16]
  assign io_arr_out_73 = arr_73; // @[fill.scala 23:16]
  assign io_arr_out_74 = arr_74; // @[fill.scala 23:16]
  assign io_arr_out_75 = arr_75; // @[fill.scala 23:16]
  assign io_arr_out_76 = arr_76; // @[fill.scala 23:16]
  assign io_arr_out_77 = arr_77; // @[fill.scala 23:16]
  assign io_arr_out_78 = arr_78; // @[fill.scala 23:16]
  assign io_arr_out_79 = arr_79; // @[fill.scala 23:16]
  assign io_ready = state == 3'h4; // @[fill.scala 50:23]
  always @(posedge clock) begin
    if (reset) begin // @[fill.scala 15:24]
      state <= 3'h7; // @[fill.scala 15:24]
    end else if (3'h7 == state) begin // @[fill.scala 25:19]
      if (io_valid) begin // @[fill.scala 27:25]
        state <= 3'h0;
      end
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      state <= 3'h1; // @[fill.scala 31:19]
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      state <= 3'h2; // @[fill.scala 35:19]
    end else begin
      state <= _GEN_563;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_0 <= _GEN_1;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h0 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_0 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_0 <= _GEN_1;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h0 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_0 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_0 <= _GEN_1;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_0 <= _GEN_241;
    end else begin
      arr_0 <= _GEN_402;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_1 <= _GEN_2;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h1 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_1 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_1 <= _GEN_2;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h1 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_1 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_1 <= _GEN_2;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_1 <= _GEN_242;
    end else begin
      arr_1 <= _GEN_403;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_2 <= _GEN_3;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h2 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_2 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_2 <= _GEN_3;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h2 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_2 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_2 <= _GEN_3;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_2 <= _GEN_243;
    end else begin
      arr_2 <= _GEN_404;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_3 <= _GEN_4;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h3 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_3 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_3 <= _GEN_4;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h3 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_3 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_3 <= _GEN_4;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_3 <= _GEN_244;
    end else begin
      arr_3 <= _GEN_405;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_4 <= _GEN_5;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h4 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_4 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_4 <= _GEN_5;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h4 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_4 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_4 <= _GEN_5;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_4 <= _GEN_245;
    end else begin
      arr_4 <= _GEN_406;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_5 <= _GEN_6;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h5 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_5 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_5 <= _GEN_6;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h5 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_5 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_5 <= _GEN_6;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_5 <= _GEN_246;
    end else begin
      arr_5 <= _GEN_407;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_6 <= _GEN_7;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h6 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_6 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_6 <= _GEN_7;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h6 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_6 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_6 <= _GEN_7;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_6 <= _GEN_247;
    end else begin
      arr_6 <= _GEN_408;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_7 <= _GEN_8;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h7 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_7 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_7 <= _GEN_8;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h7 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_7 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_7 <= _GEN_8;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_7 <= _GEN_248;
    end else begin
      arr_7 <= _GEN_409;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_8 <= _GEN_9;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h8 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_8 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_8 <= _GEN_9;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h8 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_8 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_8 <= _GEN_9;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_8 <= _GEN_249;
    end else begin
      arr_8 <= _GEN_410;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_9 <= _GEN_10;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h9 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_9 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_9 <= _GEN_10;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h9 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_9 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_9 <= _GEN_10;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_9 <= _GEN_250;
    end else begin
      arr_9 <= _GEN_411;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_10 <= _GEN_11;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'ha == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_10 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_10 <= _GEN_11;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'ha == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_10 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_10 <= _GEN_11;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_10 <= _GEN_251;
    end else begin
      arr_10 <= _GEN_412;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_11 <= _GEN_12;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'hb == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_11 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_11 <= _GEN_12;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'hb == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_11 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_11 <= _GEN_12;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_11 <= _GEN_252;
    end else begin
      arr_11 <= _GEN_413;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_12 <= _GEN_13;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'hc == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_12 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_12 <= _GEN_13;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'hc == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_12 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_12 <= _GEN_13;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_12 <= _GEN_253;
    end else begin
      arr_12 <= _GEN_414;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_13 <= _GEN_14;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'hd == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_13 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_13 <= _GEN_14;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'hd == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_13 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_13 <= _GEN_14;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_13 <= _GEN_254;
    end else begin
      arr_13 <= _GEN_415;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_14 <= _GEN_15;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'he == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_14 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_14 <= _GEN_15;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'he == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_14 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_14 <= _GEN_15;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_14 <= _GEN_255;
    end else begin
      arr_14 <= _GEN_416;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_15 <= _GEN_16;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'hf == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_15 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_15 <= _GEN_16;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'hf == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_15 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_15 <= _GEN_16;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_15 <= _GEN_256;
    end else begin
      arr_15 <= _GEN_417;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_16 <= _GEN_17;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h10 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_16 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_16 <= _GEN_17;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h10 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_16 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_16 <= _GEN_17;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_16 <= _GEN_257;
    end else begin
      arr_16 <= _GEN_418;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_17 <= _GEN_18;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h11 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_17 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_17 <= _GEN_18;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h11 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_17 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_17 <= _GEN_18;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_17 <= _GEN_258;
    end else begin
      arr_17 <= _GEN_419;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_18 <= _GEN_19;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h12 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_18 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_18 <= _GEN_19;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h12 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_18 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_18 <= _GEN_19;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_18 <= _GEN_259;
    end else begin
      arr_18 <= _GEN_420;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_19 <= _GEN_20;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h13 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_19 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_19 <= _GEN_20;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h13 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_19 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_19 <= _GEN_20;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_19 <= _GEN_260;
    end else begin
      arr_19 <= _GEN_421;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_20 <= _GEN_21;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h14 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_20 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_20 <= _GEN_21;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h14 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_20 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_20 <= _GEN_21;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_20 <= _GEN_261;
    end else begin
      arr_20 <= _GEN_422;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_21 <= _GEN_22;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h15 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_21 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_21 <= _GEN_22;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h15 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_21 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_21 <= _GEN_22;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_21 <= _GEN_262;
    end else begin
      arr_21 <= _GEN_423;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_22 <= _GEN_23;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h16 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_22 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_22 <= _GEN_23;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h16 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_22 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_22 <= _GEN_23;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_22 <= _GEN_263;
    end else begin
      arr_22 <= _GEN_424;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_23 <= _GEN_24;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h17 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_23 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_23 <= _GEN_24;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h17 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_23 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_23 <= _GEN_24;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_23 <= _GEN_264;
    end else begin
      arr_23 <= _GEN_425;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_24 <= _GEN_25;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h18 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_24 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_24 <= _GEN_25;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h18 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_24 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_24 <= _GEN_25;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_24 <= _GEN_265;
    end else begin
      arr_24 <= _GEN_426;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_25 <= _GEN_26;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h19 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_25 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_25 <= _GEN_26;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h19 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_25 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_25 <= _GEN_26;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_25 <= _GEN_266;
    end else begin
      arr_25 <= _GEN_427;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_26 <= _GEN_27;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h1a == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_26 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_26 <= _GEN_27;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h1a == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_26 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_26 <= _GEN_27;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_26 <= _GEN_267;
    end else begin
      arr_26 <= _GEN_428;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_27 <= _GEN_28;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h1b == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_27 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_27 <= _GEN_28;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h1b == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_27 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_27 <= _GEN_28;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_27 <= _GEN_268;
    end else begin
      arr_27 <= _GEN_429;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_28 <= _GEN_29;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h1c == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_28 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_28 <= _GEN_29;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h1c == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_28 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_28 <= _GEN_29;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_28 <= _GEN_269;
    end else begin
      arr_28 <= _GEN_430;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_29 <= _GEN_30;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h1d == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_29 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_29 <= _GEN_30;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h1d == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_29 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_29 <= _GEN_30;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_29 <= _GEN_270;
    end else begin
      arr_29 <= _GEN_431;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_30 <= _GEN_31;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h1e == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_30 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_30 <= _GEN_31;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h1e == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_30 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_30 <= _GEN_31;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_30 <= _GEN_271;
    end else begin
      arr_30 <= _GEN_432;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_31 <= _GEN_32;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h1f == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_31 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_31 <= _GEN_32;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h1f == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_31 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_31 <= _GEN_32;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_31 <= _GEN_272;
    end else begin
      arr_31 <= _GEN_433;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_32 <= _GEN_33;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h20 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_32 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_32 <= _GEN_33;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h20 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_32 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_32 <= _GEN_33;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_32 <= _GEN_273;
    end else begin
      arr_32 <= _GEN_434;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_33 <= _GEN_34;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h21 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_33 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_33 <= _GEN_34;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h21 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_33 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_33 <= _GEN_34;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_33 <= _GEN_274;
    end else begin
      arr_33 <= _GEN_435;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_34 <= _GEN_35;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h22 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_34 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_34 <= _GEN_35;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h22 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_34 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_34 <= _GEN_35;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_34 <= _GEN_275;
    end else begin
      arr_34 <= _GEN_436;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_35 <= _GEN_36;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h23 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_35 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_35 <= _GEN_36;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h23 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_35 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_35 <= _GEN_36;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_35 <= _GEN_276;
    end else begin
      arr_35 <= _GEN_437;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_36 <= _GEN_37;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h24 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_36 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_36 <= _GEN_37;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h24 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_36 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_36 <= _GEN_37;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_36 <= _GEN_277;
    end else begin
      arr_36 <= _GEN_438;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_37 <= _GEN_38;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h25 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_37 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_37 <= _GEN_38;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h25 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_37 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_37 <= _GEN_38;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_37 <= _GEN_278;
    end else begin
      arr_37 <= _GEN_439;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_38 <= _GEN_39;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h26 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_38 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_38 <= _GEN_39;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h26 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_38 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_38 <= _GEN_39;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_38 <= _GEN_279;
    end else begin
      arr_38 <= _GEN_440;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_39 <= _GEN_40;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h27 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_39 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_39 <= _GEN_40;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h27 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_39 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_39 <= _GEN_40;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_39 <= _GEN_280;
    end else begin
      arr_39 <= _GEN_441;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_40 <= _GEN_41;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h28 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_40 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_40 <= _GEN_41;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h28 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_40 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_40 <= _GEN_41;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_40 <= _GEN_281;
    end else begin
      arr_40 <= _GEN_442;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_41 <= _GEN_42;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h29 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_41 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_41 <= _GEN_42;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h29 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_41 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_41 <= _GEN_42;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_41 <= _GEN_282;
    end else begin
      arr_41 <= _GEN_443;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_42 <= _GEN_43;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h2a == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_42 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_42 <= _GEN_43;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h2a == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_42 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_42 <= _GEN_43;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_42 <= _GEN_283;
    end else begin
      arr_42 <= _GEN_444;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_43 <= _GEN_44;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h2b == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_43 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_43 <= _GEN_44;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h2b == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_43 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_43 <= _GEN_44;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_43 <= _GEN_284;
    end else begin
      arr_43 <= _GEN_445;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_44 <= _GEN_45;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h2c == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_44 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_44 <= _GEN_45;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h2c == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_44 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_44 <= _GEN_45;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_44 <= _GEN_285;
    end else begin
      arr_44 <= _GEN_446;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_45 <= _GEN_46;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h2d == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_45 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_45 <= _GEN_46;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h2d == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_45 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_45 <= _GEN_46;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_45 <= _GEN_286;
    end else begin
      arr_45 <= _GEN_447;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_46 <= _GEN_47;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h2e == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_46 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_46 <= _GEN_47;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h2e == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_46 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_46 <= _GEN_47;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_46 <= _GEN_287;
    end else begin
      arr_46 <= _GEN_448;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_47 <= _GEN_48;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h2f == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_47 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_47 <= _GEN_48;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h2f == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_47 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_47 <= _GEN_48;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_47 <= _GEN_288;
    end else begin
      arr_47 <= _GEN_449;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_48 <= _GEN_49;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h30 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_48 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_48 <= _GEN_49;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h30 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_48 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_48 <= _GEN_49;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_48 <= _GEN_289;
    end else begin
      arr_48 <= _GEN_450;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_49 <= _GEN_50;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h31 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_49 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_49 <= _GEN_50;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h31 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_49 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_49 <= _GEN_50;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_49 <= _GEN_290;
    end else begin
      arr_49 <= _GEN_451;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_50 <= _GEN_51;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h32 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_50 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_50 <= _GEN_51;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h32 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_50 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_50 <= _GEN_51;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_50 <= _GEN_291;
    end else begin
      arr_50 <= _GEN_452;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_51 <= _GEN_52;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h33 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_51 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_51 <= _GEN_52;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h33 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_51 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_51 <= _GEN_52;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_51 <= _GEN_292;
    end else begin
      arr_51 <= _GEN_453;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_52 <= _GEN_53;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h34 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_52 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_52 <= _GEN_53;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h34 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_52 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_52 <= _GEN_53;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_52 <= _GEN_293;
    end else begin
      arr_52 <= _GEN_454;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_53 <= _GEN_54;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h35 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_53 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_53 <= _GEN_54;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h35 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_53 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_53 <= _GEN_54;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_53 <= _GEN_294;
    end else begin
      arr_53 <= _GEN_455;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_54 <= _GEN_55;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h36 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_54 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_54 <= _GEN_55;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h36 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_54 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_54 <= _GEN_55;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_54 <= _GEN_295;
    end else begin
      arr_54 <= _GEN_456;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_55 <= _GEN_56;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h37 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_55 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_55 <= _GEN_56;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h37 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_55 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_55 <= _GEN_56;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_55 <= _GEN_296;
    end else begin
      arr_55 <= _GEN_457;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_56 <= _GEN_57;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h38 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_56 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_56 <= _GEN_57;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h38 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_56 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_56 <= _GEN_57;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_56 <= _GEN_297;
    end else begin
      arr_56 <= _GEN_458;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_57 <= _GEN_58;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h39 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_57 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_57 <= _GEN_58;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h39 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_57 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_57 <= _GEN_58;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_57 <= _GEN_298;
    end else begin
      arr_57 <= _GEN_459;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_58 <= _GEN_59;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h3a == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_58 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_58 <= _GEN_59;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h3a == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_58 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_58 <= _GEN_59;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_58 <= _GEN_299;
    end else begin
      arr_58 <= _GEN_460;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_59 <= _GEN_60;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h3b == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_59 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_59 <= _GEN_60;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h3b == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_59 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_59 <= _GEN_60;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_59 <= _GEN_300;
    end else begin
      arr_59 <= _GEN_461;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_60 <= _GEN_61;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h3c == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_60 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_60 <= _GEN_61;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h3c == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_60 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_60 <= _GEN_61;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_60 <= _GEN_301;
    end else begin
      arr_60 <= _GEN_462;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_61 <= _GEN_62;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h3d == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_61 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_61 <= _GEN_62;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h3d == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_61 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_61 <= _GEN_62;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_61 <= _GEN_302;
    end else begin
      arr_61 <= _GEN_463;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_62 <= _GEN_63;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h3e == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_62 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_62 <= _GEN_63;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h3e == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_62 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_62 <= _GEN_63;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_62 <= _GEN_303;
    end else begin
      arr_62 <= _GEN_464;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_63 <= _GEN_64;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h3f == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_63 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_63 <= _GEN_64;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h3f == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_63 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_63 <= _GEN_64;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_63 <= _GEN_304;
    end else begin
      arr_63 <= _GEN_465;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_64 <= _GEN_65;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h40 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_64 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_64 <= _GEN_65;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h40 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_64 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_64 <= _GEN_65;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_64 <= _GEN_305;
    end else begin
      arr_64 <= _GEN_466;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_65 <= _GEN_66;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h41 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_65 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_65 <= _GEN_66;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h41 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_65 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_65 <= _GEN_66;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_65 <= _GEN_306;
    end else begin
      arr_65 <= _GEN_467;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_66 <= _GEN_67;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h42 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_66 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_66 <= _GEN_67;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h42 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_66 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_66 <= _GEN_67;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_66 <= _GEN_307;
    end else begin
      arr_66 <= _GEN_468;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_67 <= _GEN_68;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h43 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_67 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_67 <= _GEN_68;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h43 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_67 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_67 <= _GEN_68;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_67 <= _GEN_308;
    end else begin
      arr_67 <= _GEN_469;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_68 <= _GEN_69;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h44 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_68 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_68 <= _GEN_69;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h44 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_68 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_68 <= _GEN_69;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_68 <= _GEN_309;
    end else begin
      arr_68 <= _GEN_470;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_69 <= _GEN_70;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h45 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_69 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_69 <= _GEN_70;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h45 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_69 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_69 <= _GEN_70;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_69 <= _GEN_310;
    end else begin
      arr_69 <= _GEN_471;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_70 <= _GEN_71;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h46 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_70 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_70 <= _GEN_71;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h46 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_70 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_70 <= _GEN_71;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_70 <= _GEN_311;
    end else begin
      arr_70 <= _GEN_472;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_71 <= _GEN_72;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h47 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_71 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_71 <= _GEN_72;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h47 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_71 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_71 <= _GEN_72;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_71 <= _GEN_312;
    end else begin
      arr_71 <= _GEN_473;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_72 <= _GEN_73;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h48 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_72 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_72 <= _GEN_73;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h48 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_72 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_72 <= _GEN_73;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_72 <= _GEN_313;
    end else begin
      arr_72 <= _GEN_474;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_73 <= _GEN_74;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h49 == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_73 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_73 <= _GEN_74;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h49 == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_73 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_73 <= _GEN_74;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_73 <= _GEN_314;
    end else begin
      arr_73 <= _GEN_475;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_74 <= _GEN_75;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h4a == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_74 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_74 <= _GEN_75;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h4a == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_74 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_74 <= _GEN_75;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_74 <= _GEN_315;
    end else begin
      arr_74 <= _GEN_476;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_75 <= _GEN_76;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h4b == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_75 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_75 <= _GEN_76;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h4b == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_75 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_75 <= _GEN_76;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_75 <= _GEN_316;
    end else begin
      arr_75 <= _GEN_477;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_76 <= _GEN_77;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h4c == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_76 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_76 <= _GEN_77;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h4c == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_76 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_76 <= _GEN_77;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_76 <= _GEN_317;
    end else begin
      arr_76 <= _GEN_478;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_77 <= _GEN_78;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h4d == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_77 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_77 <= _GEN_78;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h4d == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_77 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_77 <= _GEN_78;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_77 <= _GEN_318;
    end else begin
      arr_77 <= _GEN_479;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_78 <= _GEN_79;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h4e == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_78 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_78 <= _GEN_79;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h4e == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_78 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_78 <= _GEN_79;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_78 <= _GEN_319;
    end else begin
      arr_78 <= _GEN_480;
    end
    if (3'h7 == state) begin // @[fill.scala 25:19]
      arr_79 <= _GEN_80;
    end else if (3'h0 == state) begin // @[fill.scala 25:19]
      if (7'h4f == _T_4[6:0]) begin // @[fill.scala 30:36]
        arr_79 <= _arr_T_6; // @[fill.scala 30:36]
      end else begin
        arr_79 <= _GEN_80;
      end
    end else if (3'h1 == state) begin // @[fill.scala 25:19]
      if (7'h4f == _T_10[6:0]) begin // @[fill.scala 34:49]
        arr_79 <= _arr_T_13; // @[fill.scala 34:49]
      end else begin
        arr_79 <= _GEN_80;
      end
    end else if (3'h2 == state) begin // @[fill.scala 25:19]
      arr_79 <= _GEN_320;
    end else begin
      arr_79 <= _GEN_481;
    end
    REG <= ~io_valid; // @[fill.scala 20:18]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  arr_0 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  arr_1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  arr_2 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  arr_3 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  arr_4 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  arr_5 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  arr_6 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  arr_7 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  arr_8 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  arr_9 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  arr_10 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  arr_11 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  arr_12 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  arr_13 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  arr_14 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  arr_15 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  arr_16 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  arr_17 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  arr_18 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  arr_19 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  arr_20 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  arr_21 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  arr_22 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  arr_23 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  arr_24 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  arr_25 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  arr_26 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  arr_27 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  arr_28 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  arr_29 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  arr_30 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  arr_31 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  arr_32 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  arr_33 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  arr_34 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  arr_35 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  arr_36 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  arr_37 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  arr_38 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  arr_39 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  arr_40 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  arr_41 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  arr_42 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  arr_43 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  arr_44 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  arr_45 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  arr_46 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  arr_47 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  arr_48 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  arr_49 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  arr_50 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  arr_51 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  arr_52 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  arr_53 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  arr_54 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  arr_55 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  arr_56 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  arr_57 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  arr_58 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  arr_59 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  arr_60 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  arr_61 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  arr_62 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  arr_63 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  arr_64 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  arr_65 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  arr_66 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  arr_67 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  arr_68 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  arr_69 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  arr_70 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  arr_71 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  arr_72 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  arr_73 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  arr_74 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  arr_75 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  arr_76 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  arr_77 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  arr_78 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  arr_79 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  REG = _RAND_81[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module digest(
  input         clock,
  input         reset,
  input  [31:0] io_bytes_0,
  input  [31:0] io_bytes_1,
  input  [31:0] io_bytes_2,
  input  [31:0] io_bytes_3,
  input  [31:0] io_bytes_4,
  input  [31:0] io_bytes_5,
  input  [31:0] io_bytes_6,
  input  [31:0] io_bytes_7,
  input  [31:0] io_bytes_8,
  input  [31:0] io_bytes_9,
  input  [31:0] io_bytes_10,
  input  [31:0] io_bytes_11,
  input  [31:0] io_bytes_12,
  input  [31:0] io_bytes_13,
  input  [31:0] io_bytes_14,
  input  [31:0] io_bytes_15,
  input  [31:0] io_bytes_16,
  input  [31:0] io_bytes_17,
  input  [31:0] io_bytes_18,
  input  [31:0] io_bytes_19,
  input  [31:0] io_bytes_20,
  input  [31:0] io_bytes_21,
  input  [31:0] io_bytes_22,
  input  [31:0] io_bytes_23,
  input  [31:0] io_bytes_24,
  input  [31:0] io_bytes_25,
  input  [31:0] io_bytes_26,
  input  [31:0] io_bytes_27,
  input  [31:0] io_bytes_28,
  input  [31:0] io_bytes_29,
  input  [31:0] io_bytes_30,
  input  [31:0] io_bytes_31,
  input  [31:0] io_bytes_32,
  input  [31:0] io_bytes_33,
  input  [31:0] io_bytes_34,
  input  [31:0] io_bytes_35,
  input  [31:0] io_bytes_36,
  input  [31:0] io_bytes_37,
  input  [31:0] io_bytes_38,
  input  [31:0] io_bytes_39,
  input  [31:0] io_bytes_40,
  input  [31:0] io_bytes_41,
  input  [31:0] io_bytes_42,
  input  [31:0] io_bytes_43,
  input  [31:0] io_bytes_44,
  input  [31:0] io_bytes_45,
  input  [31:0] io_bytes_46,
  input  [31:0] io_bytes_47,
  input  [31:0] io_bytes_48,
  input  [31:0] io_bytes_49,
  input  [31:0] io_bytes_50,
  input  [31:0] io_bytes_51,
  input  [31:0] io_bytes_52,
  input  [31:0] io_bytes_53,
  input  [31:0] io_bytes_54,
  input  [31:0] io_bytes_55,
  input  [31:0] io_bytes_56,
  input  [31:0] io_bytes_57,
  input  [31:0] io_bytes_58,
  input  [31:0] io_bytes_59,
  input  [31:0] io_bytes_60,
  input  [31:0] io_bytes_61,
  input  [31:0] io_bytes_62,
  input  [31:0] io_bytes_63,
  input  [31:0] io_bytes_64,
  input  [31:0] io_bytes_65,
  input  [31:0] io_bytes_66,
  input  [31:0] io_bytes_67,
  input  [31:0] io_bytes_68,
  input  [31:0] io_bytes_69,
  input  [31:0] io_bytes_70,
  input  [31:0] io_bytes_71,
  input  [31:0] io_bytes_72,
  input  [31:0] io_bytes_73,
  input  [31:0] io_bytes_74,
  input  [31:0] io_bytes_75,
  input  [31:0] io_bytes_76,
  input  [31:0] io_bytes_77,
  input  [31:0] io_bytes_78,
  input  [31:0] io_bytes_79,
  input         io_valid,
  output [31:0] io_bytes_out_0,
  output [31:0] io_bytes_out_1,
  output [31:0] io_bytes_out_2,
  output [31:0] io_bytes_out_3,
  output [31:0] io_bytes_out_4,
  output [31:0] io_bytes_out_5,
  output [31:0] io_bytes_out_6,
  output [31:0] io_bytes_out_7,
  output [31:0] io_bytes_out_8,
  output [31:0] io_bytes_out_9,
  output [31:0] io_bytes_out_10,
  output [31:0] io_bytes_out_11,
  output [31:0] io_bytes_out_12,
  output [31:0] io_bytes_out_13,
  output [31:0] io_bytes_out_14,
  output [31:0] io_bytes_out_15,
  output [31:0] io_bytes_out_16,
  output [31:0] io_bytes_out_17,
  output [31:0] io_bytes_out_18,
  output [31:0] io_bytes_out_19,
  output [31:0] io_bytes_out_20,
  output [31:0] io_bytes_out_21,
  output [31:0] io_bytes_out_22,
  output [31:0] io_bytes_out_23,
  output [31:0] io_bytes_out_24,
  output [31:0] io_bytes_out_25,
  output [31:0] io_bytes_out_26,
  output [31:0] io_bytes_out_27,
  output [31:0] io_bytes_out_28,
  output [31:0] io_bytes_out_29,
  output [31:0] io_bytes_out_30,
  output [31:0] io_bytes_out_31,
  output [31:0] io_bytes_out_32,
  output [31:0] io_bytes_out_33,
  output [31:0] io_bytes_out_34,
  output [31:0] io_bytes_out_35,
  output [31:0] io_bytes_out_36,
  output [31:0] io_bytes_out_37,
  output [31:0] io_bytes_out_38,
  output [31:0] io_bytes_out_39,
  output [31:0] io_bytes_out_40,
  output [31:0] io_bytes_out_41,
  output [31:0] io_bytes_out_42,
  output [31:0] io_bytes_out_43,
  output [31:0] io_bytes_out_44,
  output [31:0] io_bytes_out_45,
  output [31:0] io_bytes_out_46,
  output [31:0] io_bytes_out_47,
  output [31:0] io_bytes_out_48,
  output [31:0] io_bytes_out_49,
  output [31:0] io_bytes_out_50,
  output [31:0] io_bytes_out_51,
  output [31:0] io_bytes_out_52,
  output [31:0] io_bytes_out_53,
  output [31:0] io_bytes_out_54,
  output [31:0] io_bytes_out_55,
  output [31:0] io_bytes_out_56,
  output [31:0] io_bytes_out_57,
  output [31:0] io_bytes_out_58,
  output [31:0] io_bytes_out_59,
  output [31:0] io_bytes_out_60,
  output [31:0] io_bytes_out_61,
  output [31:0] io_bytes_out_62,
  output [31:0] io_bytes_out_63,
  output [31:0] io_bytes_out_64,
  output [31:0] io_bytes_out_65,
  output [31:0] io_bytes_out_66,
  output [31:0] io_bytes_out_67,
  output [31:0] io_bytes_out_68,
  output [31:0] io_bytes_out_69,
  output [31:0] io_bytes_out_70,
  output [31:0] io_bytes_out_71,
  output [31:0] io_bytes_out_72,
  output [31:0] io_bytes_out_73,
  output [31:0] io_bytes_out_74,
  output [31:0] io_bytes_out_75,
  output [31:0] io_bytes_out_76,
  output [31:0] io_bytes_out_77,
  output [31:0] io_bytes_out_78,
  output [31:0] io_bytes_out_79,
  output        io_ready,
  output [31:0] io_out_digest_0,
  output [31:0] io_out_digest_1,
  output [31:0] io_out_digest_2,
  output [31:0] io_out_digest_3,
  output [31:0] io_out_digest_4,
  output [31:0] io_out_digest_5,
  output [31:0] io_out_digest_6,
  output [31:0] io_out_digest_7,
  output [31:0] io_out_digest_8,
  output [31:0] io_out_digest_9,
  output [31:0] io_out_digest_10,
  output [31:0] io_out_digest_11,
  output [31:0] io_out_digest_12,
  output [31:0] io_out_digest_13,
  output [31:0] io_out_digest_14,
  output [31:0] io_out_digest_15,
  output [31:0] io_out_digest_16,
  output [31:0] io_out_digest_17,
  output [31:0] io_out_digest_18,
  output [31:0] io_out_digest_19,
  output [31:0] io_out_digest_20,
  output [31:0] io_out_digest_21,
  output [31:0] io_out_digest_22,
  output [31:0] io_out_digest_23,
  output [31:0] io_out_digest_24,
  output [31:0] io_out_digest_25,
  output [31:0] io_out_digest_26,
  output [31:0] io_out_digest_27,
  output [31:0] io_out_digest_28,
  output [31:0] io_out_digest_29,
  output [31:0] io_out_digest_30,
  output [31:0] io_out_digest_31,
  output [31:0] io_out_digest_32,
  output [31:0] io_out_digest_33,
  output [31:0] io_out_digest_34,
  output [31:0] io_out_digest_35,
  output [31:0] io_out_digest_36,
  output [31:0] io_out_digest_37,
  output [31:0] io_out_digest_38,
  output [31:0] io_out_digest_39,
  output [31:0] io_out_digest_40,
  output [31:0] io_out_digest_41,
  output [31:0] io_out_digest_42,
  output [31:0] io_out_digest_43,
  output [31:0] io_out_digest_44,
  output [31:0] io_out_digest_45,
  output [31:0] io_out_digest_46,
  output [31:0] io_out_digest_47,
  output [31:0] io_out_digest_48,
  output [31:0] io_out_digest_49,
  output [31:0] io_out_digest_50,
  output [31:0] io_out_digest_51,
  output [31:0] io_out_digest_52,
  output [31:0] io_out_digest_53,
  output [31:0] io_out_digest_54,
  output [31:0] io_out_digest_55,
  output [31:0] io_out_digest_56,
  output [31:0] io_out_digest_57,
  output [31:0] io_out_digest_58,
  output [31:0] io_out_digest_59,
  output [31:0] io_out_digest_60,
  output [31:0] io_out_digest_61,
  output [31:0] io_out_digest_62,
  output [31:0] io_out_digest_63,
  output [31:0] io_out_digest_64,
  output [31:0] io_out_digest_65,
  output [31:0] io_out_digest_66,
  output [31:0] io_out_digest_67,
  output [31:0] io_out_digest_68,
  output [31:0] io_out_digest_69,
  output [31:0] io_out_digest_70,
  output [31:0] io_out_digest_71,
  output [31:0] io_out_digest_72,
  output [31:0] io_out_digest_73,
  output [31:0] io_out_digest_74,
  output [31:0] io_out_digest_75,
  output [31:0] io_out_digest_76,
  output [31:0] io_out_digest_77,
  output [31:0] io_out_digest_78,
  output [31:0] io_out_digest_79
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
`endif // RANDOMIZE_REG_INIT
  wire  __m_rol_0_clock; // @[digest.scala 41:27]
  wire  __m_rol_0_reset; // @[digest.scala 41:27]
  wire [31:0] __m_rol_0_io_num; // @[digest.scala 41:27]
  wire [31:0] __m_rol_0_io_cnt; // @[digest.scala 41:27]
  wire  __m_rol_0_io_valid; // @[digest.scala 41:27]
  wire  __m_rol_0_io_ready; // @[digest.scala 41:27]
  wire [31:0] __m_rol_0_io_out_rol; // @[digest.scala 41:27]
  wire  __m_rol_1_clock; // @[digest.scala 45:27]
  wire  __m_rol_1_reset; // @[digest.scala 45:27]
  wire [31:0] __m_rol_1_io_num; // @[digest.scala 45:27]
  wire [31:0] __m_rol_1_io_cnt; // @[digest.scala 45:27]
  wire  __m_rol_1_io_valid; // @[digest.scala 45:27]
  wire  __m_rol_1_io_ready; // @[digest.scala 45:27]
  wire [31:0] __m_rol_1_io_out_rol; // @[digest.scala 45:27]
  wire  __m_rol_2_clock; // @[digest.scala 49:27]
  wire  __m_rol_2_reset; // @[digest.scala 49:27]
  wire [31:0] __m_rol_2_io_num; // @[digest.scala 49:27]
  wire [31:0] __m_rol_2_io_cnt; // @[digest.scala 49:27]
  wire  __m_rol_2_io_valid; // @[digest.scala 49:27]
  wire  __m_rol_2_io_ready; // @[digest.scala 49:27]
  wire [31:0] __m_rol_2_io_out_rol; // @[digest.scala 49:27]
  wire  __m_fill_0_clock; // @[digest.scala 54:28]
  wire  __m_fill_0_reset; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_value; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_0; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_1; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_2; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_3; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_4; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_5; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_6; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_7; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_8; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_9; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_10; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_11; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_12; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_13; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_14; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_15; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_16; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_17; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_18; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_19; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_20; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_21; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_22; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_23; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_24; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_25; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_26; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_27; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_28; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_29; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_30; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_31; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_32; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_33; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_34; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_35; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_36; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_37; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_38; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_39; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_40; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_41; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_42; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_43; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_44; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_45; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_46; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_47; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_48; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_49; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_50; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_51; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_52; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_53; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_54; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_55; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_56; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_57; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_58; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_59; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_60; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_61; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_62; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_63; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_64; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_65; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_66; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_67; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_68; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_69; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_70; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_71; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_72; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_73; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_74; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_75; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_76; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_77; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_78; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_79; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_off; // @[digest.scala 54:28]
  wire  __m_fill_0_io_valid; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_0; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_1; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_2; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_3; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_4; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_5; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_6; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_7; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_8; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_9; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_10; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_11; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_12; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_13; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_14; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_15; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_16; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_17; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_18; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_19; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_20; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_21; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_22; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_23; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_24; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_25; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_26; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_27; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_28; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_29; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_30; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_31; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_32; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_33; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_34; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_35; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_36; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_37; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_38; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_39; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_40; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_41; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_42; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_43; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_44; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_45; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_46; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_47; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_48; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_49; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_50; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_51; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_52; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_53; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_54; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_55; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_56; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_57; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_58; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_59; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_60; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_61; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_62; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_63; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_64; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_65; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_66; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_67; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_68; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_69; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_70; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_71; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_72; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_73; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_74; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_75; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_76; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_77; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_78; // @[digest.scala 54:28]
  wire [31:0] __m_fill_0_io_arr_out_79; // @[digest.scala 54:28]
  wire  __m_fill_0_io_ready; // @[digest.scala 54:28]
  wire  __m_fill_1_clock; // @[digest.scala 59:28]
  wire  __m_fill_1_reset; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_value; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_0; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_1; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_2; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_3; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_4; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_5; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_6; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_7; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_8; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_9; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_10; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_11; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_12; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_13; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_14; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_15; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_16; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_17; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_18; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_19; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_20; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_21; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_22; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_23; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_24; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_25; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_26; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_27; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_28; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_29; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_30; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_31; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_32; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_33; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_34; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_35; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_36; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_37; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_38; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_39; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_40; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_41; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_42; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_43; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_44; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_45; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_46; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_47; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_48; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_49; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_50; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_51; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_52; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_53; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_54; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_55; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_56; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_57; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_58; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_59; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_60; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_61; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_62; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_63; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_64; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_65; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_66; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_67; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_68; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_69; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_70; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_71; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_72; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_73; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_74; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_75; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_76; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_77; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_78; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_79; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_off; // @[digest.scala 59:28]
  wire  __m_fill_1_io_valid; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_0; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_1; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_2; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_3; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_4; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_5; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_6; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_7; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_8; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_9; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_10; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_11; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_12; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_13; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_14; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_15; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_16; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_17; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_18; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_19; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_20; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_21; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_22; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_23; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_24; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_25; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_26; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_27; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_28; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_29; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_30; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_31; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_32; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_33; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_34; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_35; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_36; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_37; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_38; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_39; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_40; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_41; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_42; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_43; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_44; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_45; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_46; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_47; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_48; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_49; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_50; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_51; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_52; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_53; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_54; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_55; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_56; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_57; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_58; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_59; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_60; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_61; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_62; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_63; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_64; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_65; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_66; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_67; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_68; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_69; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_70; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_71; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_72; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_73; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_74; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_75; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_76; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_77; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_78; // @[digest.scala 59:28]
  wire [31:0] __m_fill_1_io_arr_out_79; // @[digest.scala 59:28]
  wire  __m_fill_1_io_ready; // @[digest.scala 59:28]
  wire  __m_fill_2_clock; // @[digest.scala 64:28]
  wire  __m_fill_2_reset; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_value; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_0; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_1; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_2; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_3; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_4; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_5; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_6; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_7; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_8; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_9; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_10; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_11; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_12; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_13; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_14; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_15; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_16; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_17; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_18; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_19; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_20; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_21; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_22; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_23; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_24; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_25; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_26; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_27; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_28; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_29; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_30; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_31; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_32; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_33; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_34; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_35; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_36; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_37; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_38; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_39; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_40; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_41; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_42; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_43; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_44; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_45; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_46; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_47; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_48; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_49; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_50; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_51; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_52; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_53; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_54; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_55; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_56; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_57; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_58; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_59; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_60; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_61; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_62; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_63; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_64; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_65; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_66; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_67; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_68; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_69; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_70; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_71; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_72; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_73; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_74; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_75; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_76; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_77; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_78; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_79; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_off; // @[digest.scala 64:28]
  wire  __m_fill_2_io_valid; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_0; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_1; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_2; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_3; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_4; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_5; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_6; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_7; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_8; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_9; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_10; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_11; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_12; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_13; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_14; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_15; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_16; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_17; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_18; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_19; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_20; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_21; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_22; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_23; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_24; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_25; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_26; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_27; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_28; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_29; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_30; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_31; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_32; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_33; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_34; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_35; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_36; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_37; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_38; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_39; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_40; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_41; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_42; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_43; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_44; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_45; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_46; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_47; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_48; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_49; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_50; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_51; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_52; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_53; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_54; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_55; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_56; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_57; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_58; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_59; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_60; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_61; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_62; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_63; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_64; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_65; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_66; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_67; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_68; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_69; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_70; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_71; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_72; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_73; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_74; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_75; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_76; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_77; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_78; // @[digest.scala 64:28]
  wire [31:0] __m_fill_2_io_arr_out_79; // @[digest.scala 64:28]
  wire  __m_fill_2_io_ready; // @[digest.scala 64:28]
  wire  __m_fill_3_clock; // @[digest.scala 69:28]
  wire  __m_fill_3_reset; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_value; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_0; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_1; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_2; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_3; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_4; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_5; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_6; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_7; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_8; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_9; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_10; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_11; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_12; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_13; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_14; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_15; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_16; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_17; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_18; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_19; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_20; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_21; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_22; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_23; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_24; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_25; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_26; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_27; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_28; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_29; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_30; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_31; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_32; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_33; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_34; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_35; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_36; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_37; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_38; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_39; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_40; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_41; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_42; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_43; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_44; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_45; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_46; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_47; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_48; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_49; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_50; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_51; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_52; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_53; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_54; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_55; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_56; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_57; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_58; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_59; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_60; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_61; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_62; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_63; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_64; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_65; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_66; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_67; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_68; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_69; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_70; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_71; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_72; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_73; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_74; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_75; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_76; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_77; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_78; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_79; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_off; // @[digest.scala 69:28]
  wire  __m_fill_3_io_valid; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_0; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_1; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_2; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_3; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_4; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_5; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_6; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_7; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_8; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_9; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_10; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_11; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_12; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_13; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_14; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_15; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_16; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_17; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_18; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_19; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_20; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_21; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_22; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_23; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_24; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_25; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_26; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_27; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_28; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_29; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_30; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_31; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_32; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_33; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_34; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_35; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_36; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_37; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_38; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_39; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_40; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_41; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_42; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_43; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_44; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_45; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_46; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_47; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_48; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_49; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_50; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_51; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_52; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_53; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_54; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_55; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_56; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_57; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_58; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_59; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_60; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_61; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_62; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_63; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_64; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_65; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_66; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_67; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_68; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_69; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_70; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_71; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_72; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_73; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_74; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_75; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_76; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_77; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_78; // @[digest.scala 69:28]
  wire [31:0] __m_fill_3_io_arr_out_79; // @[digest.scala 69:28]
  wire  __m_fill_3_io_ready; // @[digest.scala 69:28]
  wire  __m_fill_4_clock; // @[digest.scala 74:28]
  wire  __m_fill_4_reset; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_value; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_0; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_1; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_2; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_3; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_4; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_5; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_6; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_7; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_8; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_9; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_10; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_11; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_12; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_13; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_14; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_15; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_16; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_17; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_18; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_19; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_20; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_21; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_22; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_23; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_24; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_25; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_26; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_27; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_28; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_29; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_30; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_31; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_32; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_33; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_34; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_35; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_36; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_37; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_38; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_39; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_40; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_41; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_42; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_43; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_44; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_45; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_46; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_47; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_48; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_49; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_50; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_51; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_52; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_53; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_54; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_55; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_56; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_57; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_58; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_59; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_60; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_61; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_62; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_63; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_64; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_65; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_66; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_67; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_68; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_69; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_70; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_71; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_72; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_73; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_74; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_75; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_76; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_77; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_78; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_79; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_off; // @[digest.scala 74:28]
  wire  __m_fill_4_io_valid; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_0; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_1; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_2; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_3; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_4; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_5; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_6; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_7; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_8; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_9; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_10; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_11; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_12; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_13; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_14; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_15; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_16; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_17; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_18; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_19; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_20; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_21; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_22; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_23; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_24; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_25; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_26; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_27; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_28; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_29; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_30; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_31; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_32; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_33; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_34; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_35; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_36; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_37; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_38; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_39; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_40; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_41; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_42; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_43; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_44; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_45; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_46; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_47; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_48; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_49; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_50; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_51; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_52; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_53; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_54; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_55; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_56; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_57; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_58; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_59; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_60; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_61; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_62; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_63; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_64; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_65; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_66; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_67; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_68; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_69; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_70; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_71; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_72; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_73; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_74; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_75; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_76; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_77; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_78; // @[digest.scala 74:28]
  wire [31:0] __m_fill_4_io_arr_out_79; // @[digest.scala 74:28]
  wire  __m_fill_4_io_ready; // @[digest.scala 74:28]
  reg [5:0] state; // @[digest.scala 14:24]
  wire [5:0] _GEN_0 = reset ? 6'h3f : state; // @[digest.scala 15:26 16:15 14:24]
  reg [31:0] bytes_0; // @[digest.scala 18:20]
  reg [31:0] bytes_1; // @[digest.scala 18:20]
  reg [31:0] bytes_2; // @[digest.scala 18:20]
  reg [31:0] bytes_3; // @[digest.scala 18:20]
  reg [31:0] bytes_4; // @[digest.scala 18:20]
  reg [31:0] bytes_5; // @[digest.scala 18:20]
  reg [31:0] bytes_6; // @[digest.scala 18:20]
  reg [31:0] bytes_7; // @[digest.scala 18:20]
  reg [31:0] bytes_8; // @[digest.scala 18:20]
  reg [31:0] bytes_9; // @[digest.scala 18:20]
  reg [31:0] bytes_10; // @[digest.scala 18:20]
  reg [31:0] bytes_11; // @[digest.scala 18:20]
  reg [31:0] bytes_12; // @[digest.scala 18:20]
  reg [31:0] bytes_13; // @[digest.scala 18:20]
  reg [31:0] bytes_14; // @[digest.scala 18:20]
  reg [31:0] bytes_15; // @[digest.scala 18:20]
  reg [31:0] bytes_16; // @[digest.scala 18:20]
  reg [31:0] bytes_17; // @[digest.scala 18:20]
  reg [31:0] bytes_18; // @[digest.scala 18:20]
  reg [31:0] bytes_19; // @[digest.scala 18:20]
  reg [31:0] bytes_20; // @[digest.scala 18:20]
  reg [31:0] bytes_21; // @[digest.scala 18:20]
  reg [31:0] bytes_22; // @[digest.scala 18:20]
  reg [31:0] bytes_23; // @[digest.scala 18:20]
  reg [31:0] bytes_24; // @[digest.scala 18:20]
  reg [31:0] bytes_25; // @[digest.scala 18:20]
  reg [31:0] bytes_26; // @[digest.scala 18:20]
  reg [31:0] bytes_27; // @[digest.scala 18:20]
  reg [31:0] bytes_28; // @[digest.scala 18:20]
  reg [31:0] bytes_29; // @[digest.scala 18:20]
  reg [31:0] bytes_30; // @[digest.scala 18:20]
  reg [31:0] bytes_31; // @[digest.scala 18:20]
  reg [31:0] bytes_32; // @[digest.scala 18:20]
  reg [31:0] bytes_33; // @[digest.scala 18:20]
  reg [31:0] bytes_34; // @[digest.scala 18:20]
  reg [31:0] bytes_35; // @[digest.scala 18:20]
  reg [31:0] bytes_36; // @[digest.scala 18:20]
  reg [31:0] bytes_37; // @[digest.scala 18:20]
  reg [31:0] bytes_38; // @[digest.scala 18:20]
  reg [31:0] bytes_39; // @[digest.scala 18:20]
  reg [31:0] bytes_40; // @[digest.scala 18:20]
  reg [31:0] bytes_41; // @[digest.scala 18:20]
  reg [31:0] bytes_42; // @[digest.scala 18:20]
  reg [31:0] bytes_43; // @[digest.scala 18:20]
  reg [31:0] bytes_44; // @[digest.scala 18:20]
  reg [31:0] bytes_45; // @[digest.scala 18:20]
  reg [31:0] bytes_46; // @[digest.scala 18:20]
  reg [31:0] bytes_47; // @[digest.scala 18:20]
  reg [31:0] bytes_48; // @[digest.scala 18:20]
  reg [31:0] bytes_49; // @[digest.scala 18:20]
  reg [31:0] bytes_50; // @[digest.scala 18:20]
  reg [31:0] bytes_51; // @[digest.scala 18:20]
  reg [31:0] bytes_52; // @[digest.scala 18:20]
  reg [31:0] bytes_53; // @[digest.scala 18:20]
  reg [31:0] bytes_54; // @[digest.scala 18:20]
  reg [31:0] bytes_55; // @[digest.scala 18:20]
  reg [31:0] bytes_56; // @[digest.scala 18:20]
  reg [31:0] bytes_57; // @[digest.scala 18:20]
  reg [31:0] bytes_58; // @[digest.scala 18:20]
  reg [31:0] bytes_59; // @[digest.scala 18:20]
  reg [31:0] bytes_60; // @[digest.scala 18:20]
  reg [31:0] bytes_61; // @[digest.scala 18:20]
  reg [31:0] bytes_62; // @[digest.scala 18:20]
  reg [31:0] bytes_63; // @[digest.scala 18:20]
  reg [31:0] bytes_64; // @[digest.scala 18:20]
  reg [31:0] bytes_65; // @[digest.scala 18:20]
  reg [31:0] bytes_66; // @[digest.scala 18:20]
  reg [31:0] bytes_67; // @[digest.scala 18:20]
  reg [31:0] bytes_68; // @[digest.scala 18:20]
  reg [31:0] bytes_69; // @[digest.scala 18:20]
  reg [31:0] bytes_70; // @[digest.scala 18:20]
  reg [31:0] bytes_71; // @[digest.scala 18:20]
  reg [31:0] bytes_72; // @[digest.scala 18:20]
  reg [31:0] bytes_73; // @[digest.scala 18:20]
  reg [31:0] bytes_74; // @[digest.scala 18:20]
  reg [31:0] bytes_75; // @[digest.scala 18:20]
  reg [31:0] bytes_76; // @[digest.scala 18:20]
  reg [31:0] bytes_77; // @[digest.scala 18:20]
  reg [31:0] bytes_78; // @[digest.scala 18:20]
  reg [31:0] bytes_79; // @[digest.scala 18:20]
  reg  REG; // @[digest.scala 19:17]
  reg [31:0] i; // @[digest.scala 23:16]
  reg [31:0] a; // @[digest.scala 24:16]
  reg [31:0] b; // @[digest.scala 25:16]
  reg [31:0] c; // @[digest.scala 26:16]
  reg [31:0] d; // @[digest.scala 27:16]
  reg [31:0] e; // @[digest.scala 28:16]
  reg [31:0] olda; // @[digest.scala 29:19]
  reg [31:0] oldb; // @[digest.scala 30:19]
  reg [31:0] oldc; // @[digest.scala 31:19]
  reg [31:0] oldd; // @[digest.scala 32:19]
  reg [31:0] olde; // @[digest.scala 33:19]
  reg [31:0] j; // @[digest.scala 34:16]
  reg [31:0] t; // @[digest.scala 35:16]
  reg [31:0] blksLength; // @[digest.scala 37:25]
  reg [31:0] temp; // @[digest.scala 38:19]
  reg [31:0] blks_0; // @[digest.scala 39:19]
  reg [31:0] blks_1; // @[digest.scala 39:19]
  reg [31:0] blks_2; // @[digest.scala 39:19]
  reg [31:0] blks_3; // @[digest.scala 39:19]
  reg [31:0] blks_4; // @[digest.scala 39:19]
  reg [31:0] blks_5; // @[digest.scala 39:19]
  reg [31:0] blks_6; // @[digest.scala 39:19]
  reg [31:0] blks_7; // @[digest.scala 39:19]
  reg [31:0] blks_8; // @[digest.scala 39:19]
  reg [31:0] blks_9; // @[digest.scala 39:19]
  reg [31:0] blks_10; // @[digest.scala 39:19]
  reg [31:0] blks_11; // @[digest.scala 39:19]
  reg [31:0] blks_12; // @[digest.scala 39:19]
  reg [31:0] blks_13; // @[digest.scala 39:19]
  reg [31:0] blks_14; // @[digest.scala 39:19]
  reg [31:0] blks_15; // @[digest.scala 39:19]
  reg [31:0] blks_16; // @[digest.scala 39:19]
  reg [31:0] blks_17; // @[digest.scala 39:19]
  reg [31:0] blks_18; // @[digest.scala 39:19]
  reg [31:0] blks_19; // @[digest.scala 39:19]
  reg [31:0] blks_20; // @[digest.scala 39:19]
  reg [31:0] blks_21; // @[digest.scala 39:19]
  reg [31:0] blks_22; // @[digest.scala 39:19]
  reg [31:0] blks_23; // @[digest.scala 39:19]
  reg [31:0] blks_24; // @[digest.scala 39:19]
  reg [31:0] blks_25; // @[digest.scala 39:19]
  reg [31:0] blks_26; // @[digest.scala 39:19]
  reg [31:0] blks_27; // @[digest.scala 39:19]
  reg [31:0] blks_28; // @[digest.scala 39:19]
  reg [31:0] blks_29; // @[digest.scala 39:19]
  reg [31:0] blks_30; // @[digest.scala 39:19]
  reg [31:0] blks_31; // @[digest.scala 39:19]
  reg [31:0] blks_32; // @[digest.scala 39:19]
  reg [31:0] blks_33; // @[digest.scala 39:19]
  reg [31:0] blks_34; // @[digest.scala 39:19]
  reg [31:0] blks_35; // @[digest.scala 39:19]
  reg [31:0] blks_36; // @[digest.scala 39:19]
  reg [31:0] blks_37; // @[digest.scala 39:19]
  reg [31:0] blks_38; // @[digest.scala 39:19]
  reg [31:0] blks_39; // @[digest.scala 39:19]
  reg [31:0] blks_40; // @[digest.scala 39:19]
  reg [31:0] blks_41; // @[digest.scala 39:19]
  reg [31:0] blks_42; // @[digest.scala 39:19]
  reg [31:0] blks_43; // @[digest.scala 39:19]
  reg [31:0] blks_44; // @[digest.scala 39:19]
  reg [31:0] blks_45; // @[digest.scala 39:19]
  reg [31:0] blks_46; // @[digest.scala 39:19]
  reg [31:0] blks_47; // @[digest.scala 39:19]
  reg [31:0] blks_48; // @[digest.scala 39:19]
  reg [31:0] blks_49; // @[digest.scala 39:19]
  reg [31:0] blks_50; // @[digest.scala 39:19]
  reg [31:0] blks_51; // @[digest.scala 39:19]
  reg [31:0] blks_52; // @[digest.scala 39:19]
  reg [31:0] blks_53; // @[digest.scala 39:19]
  reg [31:0] blks_54; // @[digest.scala 39:19]
  reg [31:0] blks_55; // @[digest.scala 39:19]
  reg [31:0] blks_56; // @[digest.scala 39:19]
  reg [31:0] blks_57; // @[digest.scala 39:19]
  reg [31:0] blks_58; // @[digest.scala 39:19]
  reg [31:0] blks_59; // @[digest.scala 39:19]
  reg [31:0] blks_60; // @[digest.scala 39:19]
  reg [31:0] blks_61; // @[digest.scala 39:19]
  reg [31:0] blks_62; // @[digest.scala 39:19]
  reg [31:0] blks_63; // @[digest.scala 39:19]
  reg [31:0] blks_64; // @[digest.scala 39:19]
  reg [31:0] blks_65; // @[digest.scala 39:19]
  reg [31:0] blks_66; // @[digest.scala 39:19]
  reg [31:0] blks_67; // @[digest.scala 39:19]
  reg [31:0] blks_68; // @[digest.scala 39:19]
  reg [31:0] blks_69; // @[digest.scala 39:19]
  reg [31:0] blks_70; // @[digest.scala 39:19]
  reg [31:0] blks_71; // @[digest.scala 39:19]
  reg [31:0] blks_72; // @[digest.scala 39:19]
  reg [31:0] blks_73; // @[digest.scala 39:19]
  reg [31:0] blks_74; // @[digest.scala 39:19]
  reg [31:0] blks_75; // @[digest.scala 39:19]
  reg [31:0] blks_76; // @[digest.scala 39:19]
  reg [31:0] blks_77; // @[digest.scala 39:19]
  reg [31:0] blks_78; // @[digest.scala 39:19]
  reg [31:0] blks_79; // @[digest.scala 39:19]
  reg [31:0] w_0; // @[digest.scala 40:16]
  reg [31:0] w_1; // @[digest.scala 40:16]
  reg [31:0] w_2; // @[digest.scala 40:16]
  reg [31:0] w_3; // @[digest.scala 40:16]
  reg [31:0] w_4; // @[digest.scala 40:16]
  reg [31:0] w_5; // @[digest.scala 40:16]
  reg [31:0] w_6; // @[digest.scala 40:16]
  reg [31:0] w_7; // @[digest.scala 40:16]
  reg [31:0] w_8; // @[digest.scala 40:16]
  reg [31:0] w_9; // @[digest.scala 40:16]
  reg [31:0] w_10; // @[digest.scala 40:16]
  reg [31:0] w_11; // @[digest.scala 40:16]
  reg [31:0] w_12; // @[digest.scala 40:16]
  reg [31:0] w_13; // @[digest.scala 40:16]
  reg [31:0] w_14; // @[digest.scala 40:16]
  reg [31:0] w_15; // @[digest.scala 40:16]
  reg [31:0] w_16; // @[digest.scala 40:16]
  reg [31:0] w_17; // @[digest.scala 40:16]
  reg [31:0] w_18; // @[digest.scala 40:16]
  reg [31:0] w_19; // @[digest.scala 40:16]
  reg [31:0] w_20; // @[digest.scala 40:16]
  reg [31:0] w_21; // @[digest.scala 40:16]
  reg [31:0] w_22; // @[digest.scala 40:16]
  reg [31:0] w_23; // @[digest.scala 40:16]
  reg [31:0] w_24; // @[digest.scala 40:16]
  reg [31:0] w_25; // @[digest.scala 40:16]
  reg [31:0] w_26; // @[digest.scala 40:16]
  reg [31:0] w_27; // @[digest.scala 40:16]
  reg [31:0] w_28; // @[digest.scala 40:16]
  reg [31:0] w_29; // @[digest.scala 40:16]
  reg [31:0] w_30; // @[digest.scala 40:16]
  reg [31:0] w_31; // @[digest.scala 40:16]
  reg [31:0] w_32; // @[digest.scala 40:16]
  reg [31:0] w_33; // @[digest.scala 40:16]
  reg [31:0] w_34; // @[digest.scala 40:16]
  reg [31:0] w_35; // @[digest.scala 40:16]
  reg [31:0] w_36; // @[digest.scala 40:16]
  reg [31:0] w_37; // @[digest.scala 40:16]
  reg [31:0] w_38; // @[digest.scala 40:16]
  reg [31:0] w_39; // @[digest.scala 40:16]
  reg [31:0] w_40; // @[digest.scala 40:16]
  reg [31:0] w_41; // @[digest.scala 40:16]
  reg [31:0] w_42; // @[digest.scala 40:16]
  reg [31:0] w_43; // @[digest.scala 40:16]
  reg [31:0] w_44; // @[digest.scala 40:16]
  reg [31:0] w_45; // @[digest.scala 40:16]
  reg [31:0] w_46; // @[digest.scala 40:16]
  reg [31:0] w_47; // @[digest.scala 40:16]
  reg [31:0] w_48; // @[digest.scala 40:16]
  reg [31:0] w_49; // @[digest.scala 40:16]
  reg [31:0] w_50; // @[digest.scala 40:16]
  reg [31:0] w_51; // @[digest.scala 40:16]
  reg [31:0] w_52; // @[digest.scala 40:16]
  reg [31:0] w_53; // @[digest.scala 40:16]
  reg [31:0] w_54; // @[digest.scala 40:16]
  reg [31:0] w_55; // @[digest.scala 40:16]
  reg [31:0] w_56; // @[digest.scala 40:16]
  reg [31:0] w_57; // @[digest.scala 40:16]
  reg [31:0] w_58; // @[digest.scala 40:16]
  reg [31:0] w_59; // @[digest.scala 40:16]
  reg [31:0] w_60; // @[digest.scala 40:16]
  reg [31:0] w_61; // @[digest.scala 40:16]
  reg [31:0] w_62; // @[digest.scala 40:16]
  reg [31:0] w_63; // @[digest.scala 40:16]
  reg [31:0] w_64; // @[digest.scala 40:16]
  reg [31:0] w_65; // @[digest.scala 40:16]
  reg [31:0] w_66; // @[digest.scala 40:16]
  reg [31:0] w_67; // @[digest.scala 40:16]
  reg [31:0] w_68; // @[digest.scala 40:16]
  reg [31:0] w_69; // @[digest.scala 40:16]
  reg [31:0] w_70; // @[digest.scala 40:16]
  reg [31:0] w_71; // @[digest.scala 40:16]
  reg [31:0] w_72; // @[digest.scala 40:16]
  reg [31:0] w_73; // @[digest.scala 40:16]
  reg [31:0] w_74; // @[digest.scala 40:16]
  reg [31:0] w_75; // @[digest.scala 40:16]
  reg [31:0] w_76; // @[digest.scala 40:16]
  reg [31:0] w_77; // @[digest.scala 40:16]
  reg [31:0] w_78; // @[digest.scala 40:16]
  reg [31:0] w_79; // @[digest.scala 40:16]
  reg [31:0] digest_0; // @[digest.scala 53:21]
  reg [31:0] digest_1; // @[digest.scala 53:21]
  reg [31:0] digest_2; // @[digest.scala 53:21]
  reg [31:0] digest_3; // @[digest.scala 53:21]
  reg [31:0] digest_4; // @[digest.scala 53:21]
  reg [31:0] digest_5; // @[digest.scala 53:21]
  reg [31:0] digest_6; // @[digest.scala 53:21]
  reg [31:0] digest_7; // @[digest.scala 53:21]
  reg [31:0] digest_8; // @[digest.scala 53:21]
  reg [31:0] digest_9; // @[digest.scala 53:21]
  reg [31:0] digest_10; // @[digest.scala 53:21]
  reg [31:0] digest_11; // @[digest.scala 53:21]
  reg [31:0] digest_12; // @[digest.scala 53:21]
  reg [31:0] digest_13; // @[digest.scala 53:21]
  reg [31:0] digest_14; // @[digest.scala 53:21]
  reg [31:0] digest_15; // @[digest.scala 53:21]
  reg [31:0] digest_16; // @[digest.scala 53:21]
  reg [31:0] digest_17; // @[digest.scala 53:21]
  reg [31:0] digest_18; // @[digest.scala 53:21]
  reg [31:0] digest_19; // @[digest.scala 53:21]
  reg [31:0] digest_20; // @[digest.scala 53:21]
  reg [31:0] digest_21; // @[digest.scala 53:21]
  reg [31:0] digest_22; // @[digest.scala 53:21]
  reg [31:0] digest_23; // @[digest.scala 53:21]
  reg [31:0] digest_24; // @[digest.scala 53:21]
  reg [31:0] digest_25; // @[digest.scala 53:21]
  reg [31:0] digest_26; // @[digest.scala 53:21]
  reg [31:0] digest_27; // @[digest.scala 53:21]
  reg [31:0] digest_28; // @[digest.scala 53:21]
  reg [31:0] digest_29; // @[digest.scala 53:21]
  reg [31:0] digest_30; // @[digest.scala 53:21]
  reg [31:0] digest_31; // @[digest.scala 53:21]
  reg [31:0] digest_32; // @[digest.scala 53:21]
  reg [31:0] digest_33; // @[digest.scala 53:21]
  reg [31:0] digest_34; // @[digest.scala 53:21]
  reg [31:0] digest_35; // @[digest.scala 53:21]
  reg [31:0] digest_36; // @[digest.scala 53:21]
  reg [31:0] digest_37; // @[digest.scala 53:21]
  reg [31:0] digest_38; // @[digest.scala 53:21]
  reg [31:0] digest_39; // @[digest.scala 53:21]
  reg [31:0] digest_40; // @[digest.scala 53:21]
  reg [31:0] digest_41; // @[digest.scala 53:21]
  reg [31:0] digest_42; // @[digest.scala 53:21]
  reg [31:0] digest_43; // @[digest.scala 53:21]
  reg [31:0] digest_44; // @[digest.scala 53:21]
  reg [31:0] digest_45; // @[digest.scala 53:21]
  reg [31:0] digest_46; // @[digest.scala 53:21]
  reg [31:0] digest_47; // @[digest.scala 53:21]
  reg [31:0] digest_48; // @[digest.scala 53:21]
  reg [31:0] digest_49; // @[digest.scala 53:21]
  reg [31:0] digest_50; // @[digest.scala 53:21]
  reg [31:0] digest_51; // @[digest.scala 53:21]
  reg [31:0] digest_52; // @[digest.scala 53:21]
  reg [31:0] digest_53; // @[digest.scala 53:21]
  reg [31:0] digest_54; // @[digest.scala 53:21]
  reg [31:0] digest_55; // @[digest.scala 53:21]
  reg [31:0] digest_56; // @[digest.scala 53:21]
  reg [31:0] digest_57; // @[digest.scala 53:21]
  reg [31:0] digest_58; // @[digest.scala 53:21]
  reg [31:0] digest_59; // @[digest.scala 53:21]
  reg [31:0] digest_60; // @[digest.scala 53:21]
  reg [31:0] digest_61; // @[digest.scala 53:21]
  reg [31:0] digest_62; // @[digest.scala 53:21]
  reg [31:0] digest_63; // @[digest.scala 53:21]
  reg [31:0] digest_64; // @[digest.scala 53:21]
  reg [31:0] digest_65; // @[digest.scala 53:21]
  reg [31:0] digest_66; // @[digest.scala 53:21]
  reg [31:0] digest_67; // @[digest.scala 53:21]
  reg [31:0] digest_68; // @[digest.scala 53:21]
  reg [31:0] digest_69; // @[digest.scala 53:21]
  reg [31:0] digest_70; // @[digest.scala 53:21]
  reg [31:0] digest_71; // @[digest.scala 53:21]
  reg [31:0] digest_72; // @[digest.scala 53:21]
  reg [31:0] digest_73; // @[digest.scala 53:21]
  reg [31:0] digest_74; // @[digest.scala 53:21]
  reg [31:0] digest_75; // @[digest.scala 53:21]
  reg [31:0] digest_76; // @[digest.scala 53:21]
  reg [31:0] digest_77; // @[digest.scala 53:21]
  reg [31:0] digest_78; // @[digest.scala 53:21]
  reg [31:0] digest_79; // @[digest.scala 53:21]
  wire [63:0] _blksLength_T_6 = 32'sh1 * 32'sh10; // @[digest.scala 90:106]
  wire [64:0] _blksLength_T_7 = {{1{_blksLength_T_6[63]}},_blksLength_T_6}; // @[digest.scala 90:93]
  wire [63:0] _blksLength_T_9 = _blksLength_T_7[63:0]; // @[digest.scala 90:93]
  wire [2:0] _state_T_2 = $signed(i) < 32'sh3 ? 3'h4 : 3'h7; // @[digest.scala 98:25]
  wire [31:0] _temp_T = i; // @[digest.scala 101:38]
  wire [31:0] _temp_T_2 = $signed(i) % 32'sh4; // @[digest.scala 101:62]
  wire [63:0] _temp_T_3 = $signed(_temp_T_2) * 32'sh8; // @[digest.scala 101:75]
  wire [63:0] _temp_T_7 = 64'sh18 - $signed(_temp_T_3); // @[digest.scala 101:95]
  wire [31:0] _GEN_82 = 7'h1 == _temp_T[6:0] ? $signed(bytes_1) : $signed(bytes_0); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_83 = 7'h2 == _temp_T[6:0] ? $signed(bytes_2) : $signed(_GEN_82); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_84 = 7'h3 == _temp_T[6:0] ? $signed(bytes_3) : $signed(_GEN_83); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_85 = 7'h4 == _temp_T[6:0] ? $signed(bytes_4) : $signed(_GEN_84); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_86 = 7'h5 == _temp_T[6:0] ? $signed(bytes_5) : $signed(_GEN_85); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_87 = 7'h6 == _temp_T[6:0] ? $signed(bytes_6) : $signed(_GEN_86); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_88 = 7'h7 == _temp_T[6:0] ? $signed(bytes_7) : $signed(_GEN_87); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_89 = 7'h8 == _temp_T[6:0] ? $signed(bytes_8) : $signed(_GEN_88); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_90 = 7'h9 == _temp_T[6:0] ? $signed(bytes_9) : $signed(_GEN_89); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_91 = 7'ha == _temp_T[6:0] ? $signed(bytes_10) : $signed(_GEN_90); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_92 = 7'hb == _temp_T[6:0] ? $signed(bytes_11) : $signed(_GEN_91); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_93 = 7'hc == _temp_T[6:0] ? $signed(bytes_12) : $signed(_GEN_92); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_94 = 7'hd == _temp_T[6:0] ? $signed(bytes_13) : $signed(_GEN_93); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_95 = 7'he == _temp_T[6:0] ? $signed(bytes_14) : $signed(_GEN_94); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_96 = 7'hf == _temp_T[6:0] ? $signed(bytes_15) : $signed(_GEN_95); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_97 = 7'h10 == _temp_T[6:0] ? $signed(bytes_16) : $signed(_GEN_96); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_98 = 7'h11 == _temp_T[6:0] ? $signed(bytes_17) : $signed(_GEN_97); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_99 = 7'h12 == _temp_T[6:0] ? $signed(bytes_18) : $signed(_GEN_98); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_100 = 7'h13 == _temp_T[6:0] ? $signed(bytes_19) : $signed(_GEN_99); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_101 = 7'h14 == _temp_T[6:0] ? $signed(bytes_20) : $signed(_GEN_100); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_102 = 7'h15 == _temp_T[6:0] ? $signed(bytes_21) : $signed(_GEN_101); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_103 = 7'h16 == _temp_T[6:0] ? $signed(bytes_22) : $signed(_GEN_102); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_104 = 7'h17 == _temp_T[6:0] ? $signed(bytes_23) : $signed(_GEN_103); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_105 = 7'h18 == _temp_T[6:0] ? $signed(bytes_24) : $signed(_GEN_104); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_106 = 7'h19 == _temp_T[6:0] ? $signed(bytes_25) : $signed(_GEN_105); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_107 = 7'h1a == _temp_T[6:0] ? $signed(bytes_26) : $signed(_GEN_106); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_108 = 7'h1b == _temp_T[6:0] ? $signed(bytes_27) : $signed(_GEN_107); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_109 = 7'h1c == _temp_T[6:0] ? $signed(bytes_28) : $signed(_GEN_108); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_110 = 7'h1d == _temp_T[6:0] ? $signed(bytes_29) : $signed(_GEN_109); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_111 = 7'h1e == _temp_T[6:0] ? $signed(bytes_30) : $signed(_GEN_110); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_112 = 7'h1f == _temp_T[6:0] ? $signed(bytes_31) : $signed(_GEN_111); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_113 = 7'h20 == _temp_T[6:0] ? $signed(bytes_32) : $signed(_GEN_112); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_114 = 7'h21 == _temp_T[6:0] ? $signed(bytes_33) : $signed(_GEN_113); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_115 = 7'h22 == _temp_T[6:0] ? $signed(bytes_34) : $signed(_GEN_114); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_116 = 7'h23 == _temp_T[6:0] ? $signed(bytes_35) : $signed(_GEN_115); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_117 = 7'h24 == _temp_T[6:0] ? $signed(bytes_36) : $signed(_GEN_116); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_118 = 7'h25 == _temp_T[6:0] ? $signed(bytes_37) : $signed(_GEN_117); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_119 = 7'h26 == _temp_T[6:0] ? $signed(bytes_38) : $signed(_GEN_118); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_120 = 7'h27 == _temp_T[6:0] ? $signed(bytes_39) : $signed(_GEN_119); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_121 = 7'h28 == _temp_T[6:0] ? $signed(bytes_40) : $signed(_GEN_120); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_122 = 7'h29 == _temp_T[6:0] ? $signed(bytes_41) : $signed(_GEN_121); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_123 = 7'h2a == _temp_T[6:0] ? $signed(bytes_42) : $signed(_GEN_122); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_124 = 7'h2b == _temp_T[6:0] ? $signed(bytes_43) : $signed(_GEN_123); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_125 = 7'h2c == _temp_T[6:0] ? $signed(bytes_44) : $signed(_GEN_124); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_126 = 7'h2d == _temp_T[6:0] ? $signed(bytes_45) : $signed(_GEN_125); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_127 = 7'h2e == _temp_T[6:0] ? $signed(bytes_46) : $signed(_GEN_126); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_128 = 7'h2f == _temp_T[6:0] ? $signed(bytes_47) : $signed(_GEN_127); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_129 = 7'h30 == _temp_T[6:0] ? $signed(bytes_48) : $signed(_GEN_128); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_130 = 7'h31 == _temp_T[6:0] ? $signed(bytes_49) : $signed(_GEN_129); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_131 = 7'h32 == _temp_T[6:0] ? $signed(bytes_50) : $signed(_GEN_130); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_132 = 7'h33 == _temp_T[6:0] ? $signed(bytes_51) : $signed(_GEN_131); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_133 = 7'h34 == _temp_T[6:0] ? $signed(bytes_52) : $signed(_GEN_132); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_134 = 7'h35 == _temp_T[6:0] ? $signed(bytes_53) : $signed(_GEN_133); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_135 = 7'h36 == _temp_T[6:0] ? $signed(bytes_54) : $signed(_GEN_134); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_136 = 7'h37 == _temp_T[6:0] ? $signed(bytes_55) : $signed(_GEN_135); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_137 = 7'h38 == _temp_T[6:0] ? $signed(bytes_56) : $signed(_GEN_136); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_138 = 7'h39 == _temp_T[6:0] ? $signed(bytes_57) : $signed(_GEN_137); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_139 = 7'h3a == _temp_T[6:0] ? $signed(bytes_58) : $signed(_GEN_138); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_140 = 7'h3b == _temp_T[6:0] ? $signed(bytes_59) : $signed(_GEN_139); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_141 = 7'h3c == _temp_T[6:0] ? $signed(bytes_60) : $signed(_GEN_140); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_142 = 7'h3d == _temp_T[6:0] ? $signed(bytes_61) : $signed(_GEN_141); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_143 = 7'h3e == _temp_T[6:0] ? $signed(bytes_62) : $signed(_GEN_142); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_144 = 7'h3f == _temp_T[6:0] ? $signed(bytes_63) : $signed(_GEN_143); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_145 = 7'h40 == _temp_T[6:0] ? $signed(bytes_64) : $signed(_GEN_144); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_146 = 7'h41 == _temp_T[6:0] ? $signed(bytes_65) : $signed(_GEN_145); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_147 = 7'h42 == _temp_T[6:0] ? $signed(bytes_66) : $signed(_GEN_146); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_148 = 7'h43 == _temp_T[6:0] ? $signed(bytes_67) : $signed(_GEN_147); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_149 = 7'h44 == _temp_T[6:0] ? $signed(bytes_68) : $signed(_GEN_148); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_150 = 7'h45 == _temp_T[6:0] ? $signed(bytes_69) : $signed(_GEN_149); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_151 = 7'h46 == _temp_T[6:0] ? $signed(bytes_70) : $signed(_GEN_150); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_152 = 7'h47 == _temp_T[6:0] ? $signed(bytes_71) : $signed(_GEN_151); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_153 = 7'h48 == _temp_T[6:0] ? $signed(bytes_72) : $signed(_GEN_152); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_154 = 7'h49 == _temp_T[6:0] ? $signed(bytes_73) : $signed(_GEN_153); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_155 = 7'h4a == _temp_T[6:0] ? $signed(bytes_74) : $signed(_GEN_154); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_156 = 7'h4b == _temp_T[6:0] ? $signed(bytes_75) : $signed(_GEN_155); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_157 = 7'h4c == _temp_T[6:0] ? $signed(bytes_76) : $signed(_GEN_156); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_158 = 7'h4d == _temp_T[6:0] ? $signed(bytes_77) : $signed(_GEN_157); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_159 = 7'h4e == _temp_T[6:0] ? $signed(bytes_78) : $signed(_GEN_158); // @[digest.scala 101:{42,42}]
  wire [31:0] _GEN_160 = 7'h4f == _temp_T[6:0] ? $signed(bytes_79) : $signed(_GEN_159); // @[digest.scala 101:{42,42}]
  wire [62:0] _GEN_1 = {{31{_GEN_160[31]}},_GEN_160}; // @[digest.scala 101:42]
  wire [62:0] _temp_T_9 = $signed(_GEN_1) << _temp_T_7[4:0]; // @[digest.scala 101:42]
  wire [29:0] _GEN_34641 = i[31:2]; // @[digest.scala 105:22]
  wire [31:0] _T_12 = {{2{_GEN_34641[29]}},_GEN_34641}; // @[digest.scala 105:69]
  wire [31:0] _GEN_162 = 7'h1 == _T_12[6:0] ? $signed(blks_1) : $signed(blks_0); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_163 = 7'h2 == _T_12[6:0] ? $signed(blks_2) : $signed(_GEN_162); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_164 = 7'h3 == _T_12[6:0] ? $signed(blks_3) : $signed(_GEN_163); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_165 = 7'h4 == _T_12[6:0] ? $signed(blks_4) : $signed(_GEN_164); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_166 = 7'h5 == _T_12[6:0] ? $signed(blks_5) : $signed(_GEN_165); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_167 = 7'h6 == _T_12[6:0] ? $signed(blks_6) : $signed(_GEN_166); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_168 = 7'h7 == _T_12[6:0] ? $signed(blks_7) : $signed(_GEN_167); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_169 = 7'h8 == _T_12[6:0] ? $signed(blks_8) : $signed(_GEN_168); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_170 = 7'h9 == _T_12[6:0] ? $signed(blks_9) : $signed(_GEN_169); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_171 = 7'ha == _T_12[6:0] ? $signed(blks_10) : $signed(_GEN_170); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_172 = 7'hb == _T_12[6:0] ? $signed(blks_11) : $signed(_GEN_171); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_173 = 7'hc == _T_12[6:0] ? $signed(blks_12) : $signed(_GEN_172); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_174 = 7'hd == _T_12[6:0] ? $signed(blks_13) : $signed(_GEN_173); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_175 = 7'he == _T_12[6:0] ? $signed(blks_14) : $signed(_GEN_174); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_176 = 7'hf == _T_12[6:0] ? $signed(blks_15) : $signed(_GEN_175); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_177 = 7'h10 == _T_12[6:0] ? $signed(blks_16) : $signed(_GEN_176); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_178 = 7'h11 == _T_12[6:0] ? $signed(blks_17) : $signed(_GEN_177); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_179 = 7'h12 == _T_12[6:0] ? $signed(blks_18) : $signed(_GEN_178); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_180 = 7'h13 == _T_12[6:0] ? $signed(blks_19) : $signed(_GEN_179); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_181 = 7'h14 == _T_12[6:0] ? $signed(blks_20) : $signed(_GEN_180); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_182 = 7'h15 == _T_12[6:0] ? $signed(blks_21) : $signed(_GEN_181); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_183 = 7'h16 == _T_12[6:0] ? $signed(blks_22) : $signed(_GEN_182); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_184 = 7'h17 == _T_12[6:0] ? $signed(blks_23) : $signed(_GEN_183); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_185 = 7'h18 == _T_12[6:0] ? $signed(blks_24) : $signed(_GEN_184); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_186 = 7'h19 == _T_12[6:0] ? $signed(blks_25) : $signed(_GEN_185); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_187 = 7'h1a == _T_12[6:0] ? $signed(blks_26) : $signed(_GEN_186); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_188 = 7'h1b == _T_12[6:0] ? $signed(blks_27) : $signed(_GEN_187); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_189 = 7'h1c == _T_12[6:0] ? $signed(blks_28) : $signed(_GEN_188); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_190 = 7'h1d == _T_12[6:0] ? $signed(blks_29) : $signed(_GEN_189); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_191 = 7'h1e == _T_12[6:0] ? $signed(blks_30) : $signed(_GEN_190); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_192 = 7'h1f == _T_12[6:0] ? $signed(blks_31) : $signed(_GEN_191); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_193 = 7'h20 == _T_12[6:0] ? $signed(blks_32) : $signed(_GEN_192); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_194 = 7'h21 == _T_12[6:0] ? $signed(blks_33) : $signed(_GEN_193); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_195 = 7'h22 == _T_12[6:0] ? $signed(blks_34) : $signed(_GEN_194); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_196 = 7'h23 == _T_12[6:0] ? $signed(blks_35) : $signed(_GEN_195); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_197 = 7'h24 == _T_12[6:0] ? $signed(blks_36) : $signed(_GEN_196); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_198 = 7'h25 == _T_12[6:0] ? $signed(blks_37) : $signed(_GEN_197); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_199 = 7'h26 == _T_12[6:0] ? $signed(blks_38) : $signed(_GEN_198); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_200 = 7'h27 == _T_12[6:0] ? $signed(blks_39) : $signed(_GEN_199); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_201 = 7'h28 == _T_12[6:0] ? $signed(blks_40) : $signed(_GEN_200); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_202 = 7'h29 == _T_12[6:0] ? $signed(blks_41) : $signed(_GEN_201); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_203 = 7'h2a == _T_12[6:0] ? $signed(blks_42) : $signed(_GEN_202); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_204 = 7'h2b == _T_12[6:0] ? $signed(blks_43) : $signed(_GEN_203); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_205 = 7'h2c == _T_12[6:0] ? $signed(blks_44) : $signed(_GEN_204); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_206 = 7'h2d == _T_12[6:0] ? $signed(blks_45) : $signed(_GEN_205); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_207 = 7'h2e == _T_12[6:0] ? $signed(blks_46) : $signed(_GEN_206); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_208 = 7'h2f == _T_12[6:0] ? $signed(blks_47) : $signed(_GEN_207); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_209 = 7'h30 == _T_12[6:0] ? $signed(blks_48) : $signed(_GEN_208); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_210 = 7'h31 == _T_12[6:0] ? $signed(blks_49) : $signed(_GEN_209); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_211 = 7'h32 == _T_12[6:0] ? $signed(blks_50) : $signed(_GEN_210); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_212 = 7'h33 == _T_12[6:0] ? $signed(blks_51) : $signed(_GEN_211); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_213 = 7'h34 == _T_12[6:0] ? $signed(blks_52) : $signed(_GEN_212); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_214 = 7'h35 == _T_12[6:0] ? $signed(blks_53) : $signed(_GEN_213); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_215 = 7'h36 == _T_12[6:0] ? $signed(blks_54) : $signed(_GEN_214); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_216 = 7'h37 == _T_12[6:0] ? $signed(blks_55) : $signed(_GEN_215); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_217 = 7'h38 == _T_12[6:0] ? $signed(blks_56) : $signed(_GEN_216); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_218 = 7'h39 == _T_12[6:0] ? $signed(blks_57) : $signed(_GEN_217); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_219 = 7'h3a == _T_12[6:0] ? $signed(blks_58) : $signed(_GEN_218); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_220 = 7'h3b == _T_12[6:0] ? $signed(blks_59) : $signed(_GEN_219); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_221 = 7'h3c == _T_12[6:0] ? $signed(blks_60) : $signed(_GEN_220); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_222 = 7'h3d == _T_12[6:0] ? $signed(blks_61) : $signed(_GEN_221); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_223 = 7'h3e == _T_12[6:0] ? $signed(blks_62) : $signed(_GEN_222); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_224 = 7'h3f == _T_12[6:0] ? $signed(blks_63) : $signed(_GEN_223); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_225 = 7'h40 == _T_12[6:0] ? $signed(blks_64) : $signed(_GEN_224); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_226 = 7'h41 == _T_12[6:0] ? $signed(blks_65) : $signed(_GEN_225); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_227 = 7'h42 == _T_12[6:0] ? $signed(blks_66) : $signed(_GEN_226); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_228 = 7'h43 == _T_12[6:0] ? $signed(blks_67) : $signed(_GEN_227); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_229 = 7'h44 == _T_12[6:0] ? $signed(blks_68) : $signed(_GEN_228); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_230 = 7'h45 == _T_12[6:0] ? $signed(blks_69) : $signed(_GEN_229); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_231 = 7'h46 == _T_12[6:0] ? $signed(blks_70) : $signed(_GEN_230); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_232 = 7'h47 == _T_12[6:0] ? $signed(blks_71) : $signed(_GEN_231); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_233 = 7'h48 == _T_12[6:0] ? $signed(blks_72) : $signed(_GEN_232); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_234 = 7'h49 == _T_12[6:0] ? $signed(blks_73) : $signed(_GEN_233); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_235 = 7'h4a == _T_12[6:0] ? $signed(blks_74) : $signed(_GEN_234); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_236 = 7'h4b == _T_12[6:0] ? $signed(blks_75) : $signed(_GEN_235); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_237 = 7'h4c == _T_12[6:0] ? $signed(blks_76) : $signed(_GEN_236); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_238 = 7'h4d == _T_12[6:0] ? $signed(blks_77) : $signed(_GEN_237); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_239 = 7'h4e == _T_12[6:0] ? $signed(blks_78) : $signed(_GEN_238); // @[digest.scala 105:{136,136}]
  wire [31:0] _GEN_240 = 7'h4f == _T_12[6:0] ? $signed(blks_79) : $signed(_GEN_239); // @[digest.scala 105:{136,136}]
  wire [31:0] _blks_T_6 = $signed(_GEN_240) | $signed(temp); // @[digest.scala 105:136]
  wire [31:0] _GEN_241 = 7'h0 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_0); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_242 = 7'h1 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_1); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_243 = 7'h2 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_2); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_244 = 7'h3 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_3); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_245 = 7'h4 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_4); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_246 = 7'h5 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_5); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_247 = 7'h6 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_6); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_248 = 7'h7 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_7); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_249 = 7'h8 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_8); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_250 = 7'h9 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_9); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_251 = 7'ha == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_10); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_252 = 7'hb == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_11); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_253 = 7'hc == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_12); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_254 = 7'hd == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_13); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_255 = 7'he == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_14); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_256 = 7'hf == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_15); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_257 = 7'h10 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_16); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_258 = 7'h11 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_17); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_259 = 7'h12 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_18); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_260 = 7'h13 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_19); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_261 = 7'h14 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_20); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_262 = 7'h15 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_21); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_263 = 7'h16 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_22); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_264 = 7'h17 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_23); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_265 = 7'h18 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_24); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_266 = 7'h19 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_25); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_267 = 7'h1a == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_26); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_268 = 7'h1b == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_27); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_269 = 7'h1c == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_28); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_270 = 7'h1d == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_29); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_271 = 7'h1e == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_30); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_272 = 7'h1f == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_31); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_273 = 7'h20 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_32); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_274 = 7'h21 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_33); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_275 = 7'h22 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_34); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_276 = 7'h23 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_35); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_277 = 7'h24 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_36); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_278 = 7'h25 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_37); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_279 = 7'h26 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_38); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_280 = 7'h27 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_39); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_281 = 7'h28 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_40); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_282 = 7'h29 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_41); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_283 = 7'h2a == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_42); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_284 = 7'h2b == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_43); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_285 = 7'h2c == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_44); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_286 = 7'h2d == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_45); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_287 = 7'h2e == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_46); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_288 = 7'h2f == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_47); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_289 = 7'h30 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_48); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_290 = 7'h31 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_49); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_291 = 7'h32 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_50); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_292 = 7'h33 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_51); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_293 = 7'h34 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_52); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_294 = 7'h35 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_53); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_295 = 7'h36 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_54); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_296 = 7'h37 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_55); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_297 = 7'h38 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_56); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_298 = 7'h39 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_57); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_299 = 7'h3a == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_58); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_300 = 7'h3b == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_59); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_301 = 7'h3c == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_60); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_302 = 7'h3d == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_61); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_303 = 7'h3e == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_62); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_304 = 7'h3f == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_63); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_305 = 7'h40 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_64); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_306 = 7'h41 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_65); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_307 = 7'h42 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_66); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_308 = 7'h43 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_67); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_309 = 7'h44 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_68); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_310 = 7'h45 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_69); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_311 = 7'h46 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_70); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_312 = 7'h47 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_71); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_313 = 7'h48 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_72); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_314 = 7'h49 == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_73); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_315 = 7'h4a == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_74); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_316 = 7'h4b == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_75); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_317 = 7'h4c == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_76); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_318 = 7'h4d == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_77); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_319 = 7'h4e == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_78); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _GEN_320 = 7'h4f == _T_12[6:0] ? $signed(_blks_T_6) : $signed(blks_79); // @[digest.scala 105:{73,73} 39:19]
  wire [31:0] _i_T_2 = $signed(i) + 32'sh1; // @[digest.scala 109:21]
  wire [62:0] _temp_T_17 = 63'sh80 << _temp_T_7[4:0]; // @[digest.scala 113:35]
  wire [31:0] _T_26 = $signed(blksLength) - 32'sh1; // @[digest.scala 121:50]
  wire [63:0] _blks_T_14 = 32'sh3 * 32'sh8; // @[digest.scala 121:69]
  wire [31:0] _blks_T_27 = _blks_T_14[31:0]; // @[digest.scala 121:{54,54}]
  wire [31:0] _GEN_481 = 7'h0 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_0); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_482 = 7'h1 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_1); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_483 = 7'h2 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_2); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_484 = 7'h3 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_3); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_485 = 7'h4 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_4); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_486 = 7'h5 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_5); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_487 = 7'h6 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_6); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_488 = 7'h7 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_7); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_489 = 7'h8 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_8); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_490 = 7'h9 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_9); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_491 = 7'ha == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_10); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_492 = 7'hb == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_11); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_493 = 7'hc == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_12); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_494 = 7'hd == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_13); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_495 = 7'he == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_14); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_496 = 7'hf == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_15); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_497 = 7'h10 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_16); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_498 = 7'h11 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_17); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_499 = 7'h12 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_18); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_500 = 7'h13 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_19); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_501 = 7'h14 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_20); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_502 = 7'h15 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_21); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_503 = 7'h16 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_22); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_504 = 7'h17 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_23); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_505 = 7'h18 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_24); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_506 = 7'h19 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_25); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_507 = 7'h1a == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_26); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_508 = 7'h1b == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_27); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_509 = 7'h1c == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_28); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_510 = 7'h1d == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_29); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_511 = 7'h1e == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_30); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_512 = 7'h1f == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_31); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_513 = 7'h20 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_32); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_514 = 7'h21 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_33); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_515 = 7'h22 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_34); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_516 = 7'h23 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_35); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_517 = 7'h24 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_36); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_518 = 7'h25 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_37); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_519 = 7'h26 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_38); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_520 = 7'h27 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_39); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_521 = 7'h28 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_40); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_522 = 7'h29 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_41); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_523 = 7'h2a == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_42); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_524 = 7'h2b == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_43); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_525 = 7'h2c == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_44); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_526 = 7'h2d == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_45); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_527 = 7'h2e == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_46); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_528 = 7'h2f == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_47); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_529 = 7'h30 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_48); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_530 = 7'h31 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_49); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_531 = 7'h32 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_50); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_532 = 7'h33 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_51); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_533 = 7'h34 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_52); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_534 = 7'h35 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_53); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_535 = 7'h36 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_54); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_536 = 7'h37 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_55); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_537 = 7'h38 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_56); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_538 = 7'h39 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_57); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_539 = 7'h3a == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_58); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_540 = 7'h3b == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_59); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_541 = 7'h3c == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_60); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_542 = 7'h3d == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_61); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_543 = 7'h3e == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_62); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_544 = 7'h3f == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_63); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_545 = 7'h40 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_64); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_546 = 7'h41 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_65); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_547 = 7'h42 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_66); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_548 = 7'h43 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_67); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_549 = 7'h44 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_68); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_550 = 7'h45 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_69); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_551 = 7'h46 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_70); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_552 = 7'h47 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_71); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_553 = 7'h48 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_72); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_554 = 7'h49 == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_73); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_555 = 7'h4a == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_74); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_556 = 7'h4b == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_75); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_557 = 7'h4c == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_76); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_558 = 7'h4d == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_77); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_559 = 7'h4e == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_78); // @[digest.scala 121:{54,54} 39:19]
  wire [31:0] _GEN_560 = 7'h4f == _T_26[6:0] ? $signed(_blks_T_27) : $signed(blks_79); // @[digest.scala 121:{54,54} 39:19]
  wire [5:0] _state_T_4 = $signed(i) < $signed(blksLength) ? 6'h11 : 6'h36; // @[digest.scala 149:25]
  wire [5:0] _state_T_6 = $signed(j) < 32'sh50 ? 6'h18 : 6'h30; // @[digest.scala 176:25]
  wire [4:0] _state_T_8 = $signed(j) < 32'sh10 ? 5'h19 : 5'h1a; // @[digest.scala 179:25]
  wire [31:0] _T_44 = j; // @[digest.scala 182:25]
  wire [31:0] _w_T_3 = $signed(i) + $signed(j); // @[digest.scala 182:51]
  wire [31:0] _GEN_642 = 7'h1 == _w_T_3[6:0] ? $signed(blks_1) : $signed(blks_0); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_643 = 7'h2 == _w_T_3[6:0] ? $signed(blks_2) : $signed(_GEN_642); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_644 = 7'h3 == _w_T_3[6:0] ? $signed(blks_3) : $signed(_GEN_643); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_645 = 7'h4 == _w_T_3[6:0] ? $signed(blks_4) : $signed(_GEN_644); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_646 = 7'h5 == _w_T_3[6:0] ? $signed(blks_5) : $signed(_GEN_645); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_647 = 7'h6 == _w_T_3[6:0] ? $signed(blks_6) : $signed(_GEN_646); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_648 = 7'h7 == _w_T_3[6:0] ? $signed(blks_7) : $signed(_GEN_647); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_649 = 7'h8 == _w_T_3[6:0] ? $signed(blks_8) : $signed(_GEN_648); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_650 = 7'h9 == _w_T_3[6:0] ? $signed(blks_9) : $signed(_GEN_649); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_651 = 7'ha == _w_T_3[6:0] ? $signed(blks_10) : $signed(_GEN_650); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_652 = 7'hb == _w_T_3[6:0] ? $signed(blks_11) : $signed(_GEN_651); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_653 = 7'hc == _w_T_3[6:0] ? $signed(blks_12) : $signed(_GEN_652); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_654 = 7'hd == _w_T_3[6:0] ? $signed(blks_13) : $signed(_GEN_653); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_655 = 7'he == _w_T_3[6:0] ? $signed(blks_14) : $signed(_GEN_654); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_656 = 7'hf == _w_T_3[6:0] ? $signed(blks_15) : $signed(_GEN_655); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_657 = 7'h10 == _w_T_3[6:0] ? $signed(blks_16) : $signed(_GEN_656); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_658 = 7'h11 == _w_T_3[6:0] ? $signed(blks_17) : $signed(_GEN_657); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_659 = 7'h12 == _w_T_3[6:0] ? $signed(blks_18) : $signed(_GEN_658); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_660 = 7'h13 == _w_T_3[6:0] ? $signed(blks_19) : $signed(_GEN_659); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_661 = 7'h14 == _w_T_3[6:0] ? $signed(blks_20) : $signed(_GEN_660); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_662 = 7'h15 == _w_T_3[6:0] ? $signed(blks_21) : $signed(_GEN_661); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_663 = 7'h16 == _w_T_3[6:0] ? $signed(blks_22) : $signed(_GEN_662); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_664 = 7'h17 == _w_T_3[6:0] ? $signed(blks_23) : $signed(_GEN_663); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_665 = 7'h18 == _w_T_3[6:0] ? $signed(blks_24) : $signed(_GEN_664); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_666 = 7'h19 == _w_T_3[6:0] ? $signed(blks_25) : $signed(_GEN_665); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_667 = 7'h1a == _w_T_3[6:0] ? $signed(blks_26) : $signed(_GEN_666); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_668 = 7'h1b == _w_T_3[6:0] ? $signed(blks_27) : $signed(_GEN_667); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_669 = 7'h1c == _w_T_3[6:0] ? $signed(blks_28) : $signed(_GEN_668); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_670 = 7'h1d == _w_T_3[6:0] ? $signed(blks_29) : $signed(_GEN_669); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_671 = 7'h1e == _w_T_3[6:0] ? $signed(blks_30) : $signed(_GEN_670); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_672 = 7'h1f == _w_T_3[6:0] ? $signed(blks_31) : $signed(_GEN_671); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_673 = 7'h20 == _w_T_3[6:0] ? $signed(blks_32) : $signed(_GEN_672); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_674 = 7'h21 == _w_T_3[6:0] ? $signed(blks_33) : $signed(_GEN_673); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_675 = 7'h22 == _w_T_3[6:0] ? $signed(blks_34) : $signed(_GEN_674); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_676 = 7'h23 == _w_T_3[6:0] ? $signed(blks_35) : $signed(_GEN_675); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_677 = 7'h24 == _w_T_3[6:0] ? $signed(blks_36) : $signed(_GEN_676); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_678 = 7'h25 == _w_T_3[6:0] ? $signed(blks_37) : $signed(_GEN_677); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_679 = 7'h26 == _w_T_3[6:0] ? $signed(blks_38) : $signed(_GEN_678); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_680 = 7'h27 == _w_T_3[6:0] ? $signed(blks_39) : $signed(_GEN_679); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_681 = 7'h28 == _w_T_3[6:0] ? $signed(blks_40) : $signed(_GEN_680); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_682 = 7'h29 == _w_T_3[6:0] ? $signed(blks_41) : $signed(_GEN_681); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_683 = 7'h2a == _w_T_3[6:0] ? $signed(blks_42) : $signed(_GEN_682); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_684 = 7'h2b == _w_T_3[6:0] ? $signed(blks_43) : $signed(_GEN_683); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_685 = 7'h2c == _w_T_3[6:0] ? $signed(blks_44) : $signed(_GEN_684); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_686 = 7'h2d == _w_T_3[6:0] ? $signed(blks_45) : $signed(_GEN_685); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_687 = 7'h2e == _w_T_3[6:0] ? $signed(blks_46) : $signed(_GEN_686); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_688 = 7'h2f == _w_T_3[6:0] ? $signed(blks_47) : $signed(_GEN_687); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_689 = 7'h30 == _w_T_3[6:0] ? $signed(blks_48) : $signed(_GEN_688); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_690 = 7'h31 == _w_T_3[6:0] ? $signed(blks_49) : $signed(_GEN_689); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_691 = 7'h32 == _w_T_3[6:0] ? $signed(blks_50) : $signed(_GEN_690); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_692 = 7'h33 == _w_T_3[6:0] ? $signed(blks_51) : $signed(_GEN_691); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_693 = 7'h34 == _w_T_3[6:0] ? $signed(blks_52) : $signed(_GEN_692); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_694 = 7'h35 == _w_T_3[6:0] ? $signed(blks_53) : $signed(_GEN_693); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_695 = 7'h36 == _w_T_3[6:0] ? $signed(blks_54) : $signed(_GEN_694); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_696 = 7'h37 == _w_T_3[6:0] ? $signed(blks_55) : $signed(_GEN_695); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_697 = 7'h38 == _w_T_3[6:0] ? $signed(blks_56) : $signed(_GEN_696); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_698 = 7'h39 == _w_T_3[6:0] ? $signed(blks_57) : $signed(_GEN_697); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_699 = 7'h3a == _w_T_3[6:0] ? $signed(blks_58) : $signed(_GEN_698); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_700 = 7'h3b == _w_T_3[6:0] ? $signed(blks_59) : $signed(_GEN_699); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_701 = 7'h3c == _w_T_3[6:0] ? $signed(blks_60) : $signed(_GEN_700); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_702 = 7'h3d == _w_T_3[6:0] ? $signed(blks_61) : $signed(_GEN_701); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_703 = 7'h3e == _w_T_3[6:0] ? $signed(blks_62) : $signed(_GEN_702); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_704 = 7'h3f == _w_T_3[6:0] ? $signed(blks_63) : $signed(_GEN_703); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_705 = 7'h40 == _w_T_3[6:0] ? $signed(blks_64) : $signed(_GEN_704); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_706 = 7'h41 == _w_T_3[6:0] ? $signed(blks_65) : $signed(_GEN_705); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_707 = 7'h42 == _w_T_3[6:0] ? $signed(blks_66) : $signed(_GEN_706); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_708 = 7'h43 == _w_T_3[6:0] ? $signed(blks_67) : $signed(_GEN_707); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_709 = 7'h44 == _w_T_3[6:0] ? $signed(blks_68) : $signed(_GEN_708); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_710 = 7'h45 == _w_T_3[6:0] ? $signed(blks_69) : $signed(_GEN_709); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_711 = 7'h46 == _w_T_3[6:0] ? $signed(blks_70) : $signed(_GEN_710); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_712 = 7'h47 == _w_T_3[6:0] ? $signed(blks_71) : $signed(_GEN_711); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_713 = 7'h48 == _w_T_3[6:0] ? $signed(blks_72) : $signed(_GEN_712); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_714 = 7'h49 == _w_T_3[6:0] ? $signed(blks_73) : $signed(_GEN_713); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_715 = 7'h4a == _w_T_3[6:0] ? $signed(blks_74) : $signed(_GEN_714); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_716 = 7'h4b == _w_T_3[6:0] ? $signed(blks_75) : $signed(_GEN_715); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_717 = 7'h4c == _w_T_3[6:0] ? $signed(blks_76) : $signed(_GEN_716); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_718 = 7'h4d == _w_T_3[6:0] ? $signed(blks_77) : $signed(_GEN_717); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_719 = 7'h4e == _w_T_3[6:0] ? $signed(blks_78) : $signed(_GEN_718); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_720 = 7'h4f == _w_T_3[6:0] ? $signed(blks_79) : $signed(_GEN_719); // @[digest.scala 182:{29,29}]
  wire [31:0] _GEN_561 = 7'h0 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_0); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_562 = 7'h1 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_1); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_563 = 7'h2 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_2); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_564 = 7'h3 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_3); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_565 = 7'h4 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_4); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_566 = 7'h5 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_5); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_567 = 7'h6 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_6); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_568 = 7'h7 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_7); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_569 = 7'h8 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_8); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_570 = 7'h9 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_9); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_571 = 7'ha == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_10); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_572 = 7'hb == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_11); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_573 = 7'hc == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_12); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_574 = 7'hd == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_13); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_575 = 7'he == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_14); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_576 = 7'hf == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_15); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_577 = 7'h10 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_16); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_578 = 7'h11 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_17); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_579 = 7'h12 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_18); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_580 = 7'h13 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_19); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_581 = 7'h14 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_20); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_582 = 7'h15 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_21); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_583 = 7'h16 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_22); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_584 = 7'h17 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_23); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_585 = 7'h18 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_24); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_586 = 7'h19 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_25); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_587 = 7'h1a == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_26); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_588 = 7'h1b == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_27); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_589 = 7'h1c == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_28); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_590 = 7'h1d == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_29); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_591 = 7'h1e == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_30); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_592 = 7'h1f == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_31); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_593 = 7'h20 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_32); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_594 = 7'h21 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_33); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_595 = 7'h22 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_34); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_596 = 7'h23 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_35); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_597 = 7'h24 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_36); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_598 = 7'h25 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_37); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_599 = 7'h26 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_38); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_600 = 7'h27 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_39); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_601 = 7'h28 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_40); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_602 = 7'h29 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_41); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_603 = 7'h2a == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_42); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_604 = 7'h2b == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_43); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_605 = 7'h2c == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_44); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_606 = 7'h2d == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_45); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_607 = 7'h2e == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_46); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_608 = 7'h2f == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_47); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_609 = 7'h30 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_48); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_610 = 7'h31 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_49); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_611 = 7'h32 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_50); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_612 = 7'h33 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_51); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_613 = 7'h34 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_52); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_614 = 7'h35 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_53); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_615 = 7'h36 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_54); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_616 = 7'h37 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_55); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_617 = 7'h38 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_56); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_618 = 7'h39 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_57); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_619 = 7'h3a == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_58); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_620 = 7'h3b == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_59); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_621 = 7'h3c == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_60); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_622 = 7'h3d == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_61); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_623 = 7'h3e == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_62); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_624 = 7'h3f == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_63); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_625 = 7'h40 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_64); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_626 = 7'h41 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_65); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_627 = 7'h42 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_66); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_628 = 7'h43 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_67); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_629 = 7'h44 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_68); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_630 = 7'h45 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_69); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_631 = 7'h46 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_70); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_632 = 7'h47 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_71); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_633 = 7'h48 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_72); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_634 = 7'h49 == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_73); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_635 = 7'h4a == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_74); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_636 = 7'h4b == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_75); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_637 = 7'h4c == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_76); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_638 = 7'h4d == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_77); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_639 = 7'h4e == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_78); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _GEN_640 = 7'h4f == _T_44[6:0] ? $signed(_GEN_720) : $signed(w_79); // @[digest.scala 182:{29,29} 40:16]
  wire [31:0] _temp_T_21 = $signed(j) - 32'sh3; // @[digest.scala 186:46]
  wire [31:0] _temp_T_26 = $signed(j) - 32'sh8; // @[digest.scala 186:77]
  wire [31:0] _GEN_722 = 7'h1 == _temp_T_21[6:0] ? $signed(w_1) : $signed(w_0); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_723 = 7'h2 == _temp_T_21[6:0] ? $signed(w_2) : $signed(_GEN_722); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_724 = 7'h3 == _temp_T_21[6:0] ? $signed(w_3) : $signed(_GEN_723); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_725 = 7'h4 == _temp_T_21[6:0] ? $signed(w_4) : $signed(_GEN_724); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_726 = 7'h5 == _temp_T_21[6:0] ? $signed(w_5) : $signed(_GEN_725); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_727 = 7'h6 == _temp_T_21[6:0] ? $signed(w_6) : $signed(_GEN_726); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_728 = 7'h7 == _temp_T_21[6:0] ? $signed(w_7) : $signed(_GEN_727); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_729 = 7'h8 == _temp_T_21[6:0] ? $signed(w_8) : $signed(_GEN_728); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_730 = 7'h9 == _temp_T_21[6:0] ? $signed(w_9) : $signed(_GEN_729); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_731 = 7'ha == _temp_T_21[6:0] ? $signed(w_10) : $signed(_GEN_730); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_732 = 7'hb == _temp_T_21[6:0] ? $signed(w_11) : $signed(_GEN_731); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_733 = 7'hc == _temp_T_21[6:0] ? $signed(w_12) : $signed(_GEN_732); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_734 = 7'hd == _temp_T_21[6:0] ? $signed(w_13) : $signed(_GEN_733); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_735 = 7'he == _temp_T_21[6:0] ? $signed(w_14) : $signed(_GEN_734); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_736 = 7'hf == _temp_T_21[6:0] ? $signed(w_15) : $signed(_GEN_735); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_737 = 7'h10 == _temp_T_21[6:0] ? $signed(w_16) : $signed(_GEN_736); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_738 = 7'h11 == _temp_T_21[6:0] ? $signed(w_17) : $signed(_GEN_737); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_739 = 7'h12 == _temp_T_21[6:0] ? $signed(w_18) : $signed(_GEN_738); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_740 = 7'h13 == _temp_T_21[6:0] ? $signed(w_19) : $signed(_GEN_739); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_741 = 7'h14 == _temp_T_21[6:0] ? $signed(w_20) : $signed(_GEN_740); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_742 = 7'h15 == _temp_T_21[6:0] ? $signed(w_21) : $signed(_GEN_741); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_743 = 7'h16 == _temp_T_21[6:0] ? $signed(w_22) : $signed(_GEN_742); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_744 = 7'h17 == _temp_T_21[6:0] ? $signed(w_23) : $signed(_GEN_743); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_745 = 7'h18 == _temp_T_21[6:0] ? $signed(w_24) : $signed(_GEN_744); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_746 = 7'h19 == _temp_T_21[6:0] ? $signed(w_25) : $signed(_GEN_745); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_747 = 7'h1a == _temp_T_21[6:0] ? $signed(w_26) : $signed(_GEN_746); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_748 = 7'h1b == _temp_T_21[6:0] ? $signed(w_27) : $signed(_GEN_747); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_749 = 7'h1c == _temp_T_21[6:0] ? $signed(w_28) : $signed(_GEN_748); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_750 = 7'h1d == _temp_T_21[6:0] ? $signed(w_29) : $signed(_GEN_749); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_751 = 7'h1e == _temp_T_21[6:0] ? $signed(w_30) : $signed(_GEN_750); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_752 = 7'h1f == _temp_T_21[6:0] ? $signed(w_31) : $signed(_GEN_751); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_753 = 7'h20 == _temp_T_21[6:0] ? $signed(w_32) : $signed(_GEN_752); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_754 = 7'h21 == _temp_T_21[6:0] ? $signed(w_33) : $signed(_GEN_753); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_755 = 7'h22 == _temp_T_21[6:0] ? $signed(w_34) : $signed(_GEN_754); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_756 = 7'h23 == _temp_T_21[6:0] ? $signed(w_35) : $signed(_GEN_755); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_757 = 7'h24 == _temp_T_21[6:0] ? $signed(w_36) : $signed(_GEN_756); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_758 = 7'h25 == _temp_T_21[6:0] ? $signed(w_37) : $signed(_GEN_757); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_759 = 7'h26 == _temp_T_21[6:0] ? $signed(w_38) : $signed(_GEN_758); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_760 = 7'h27 == _temp_T_21[6:0] ? $signed(w_39) : $signed(_GEN_759); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_761 = 7'h28 == _temp_T_21[6:0] ? $signed(w_40) : $signed(_GEN_760); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_762 = 7'h29 == _temp_T_21[6:0] ? $signed(w_41) : $signed(_GEN_761); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_763 = 7'h2a == _temp_T_21[6:0] ? $signed(w_42) : $signed(_GEN_762); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_764 = 7'h2b == _temp_T_21[6:0] ? $signed(w_43) : $signed(_GEN_763); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_765 = 7'h2c == _temp_T_21[6:0] ? $signed(w_44) : $signed(_GEN_764); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_766 = 7'h2d == _temp_T_21[6:0] ? $signed(w_45) : $signed(_GEN_765); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_767 = 7'h2e == _temp_T_21[6:0] ? $signed(w_46) : $signed(_GEN_766); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_768 = 7'h2f == _temp_T_21[6:0] ? $signed(w_47) : $signed(_GEN_767); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_769 = 7'h30 == _temp_T_21[6:0] ? $signed(w_48) : $signed(_GEN_768); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_770 = 7'h31 == _temp_T_21[6:0] ? $signed(w_49) : $signed(_GEN_769); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_771 = 7'h32 == _temp_T_21[6:0] ? $signed(w_50) : $signed(_GEN_770); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_772 = 7'h33 == _temp_T_21[6:0] ? $signed(w_51) : $signed(_GEN_771); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_773 = 7'h34 == _temp_T_21[6:0] ? $signed(w_52) : $signed(_GEN_772); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_774 = 7'h35 == _temp_T_21[6:0] ? $signed(w_53) : $signed(_GEN_773); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_775 = 7'h36 == _temp_T_21[6:0] ? $signed(w_54) : $signed(_GEN_774); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_776 = 7'h37 == _temp_T_21[6:0] ? $signed(w_55) : $signed(_GEN_775); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_777 = 7'h38 == _temp_T_21[6:0] ? $signed(w_56) : $signed(_GEN_776); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_778 = 7'h39 == _temp_T_21[6:0] ? $signed(w_57) : $signed(_GEN_777); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_779 = 7'h3a == _temp_T_21[6:0] ? $signed(w_58) : $signed(_GEN_778); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_780 = 7'h3b == _temp_T_21[6:0] ? $signed(w_59) : $signed(_GEN_779); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_781 = 7'h3c == _temp_T_21[6:0] ? $signed(w_60) : $signed(_GEN_780); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_782 = 7'h3d == _temp_T_21[6:0] ? $signed(w_61) : $signed(_GEN_781); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_783 = 7'h3e == _temp_T_21[6:0] ? $signed(w_62) : $signed(_GEN_782); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_784 = 7'h3f == _temp_T_21[6:0] ? $signed(w_63) : $signed(_GEN_783); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_785 = 7'h40 == _temp_T_21[6:0] ? $signed(w_64) : $signed(_GEN_784); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_786 = 7'h41 == _temp_T_21[6:0] ? $signed(w_65) : $signed(_GEN_785); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_787 = 7'h42 == _temp_T_21[6:0] ? $signed(w_66) : $signed(_GEN_786); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_788 = 7'h43 == _temp_T_21[6:0] ? $signed(w_67) : $signed(_GEN_787); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_789 = 7'h44 == _temp_T_21[6:0] ? $signed(w_68) : $signed(_GEN_788); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_790 = 7'h45 == _temp_T_21[6:0] ? $signed(w_69) : $signed(_GEN_789); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_791 = 7'h46 == _temp_T_21[6:0] ? $signed(w_70) : $signed(_GEN_790); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_792 = 7'h47 == _temp_T_21[6:0] ? $signed(w_71) : $signed(_GEN_791); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_793 = 7'h48 == _temp_T_21[6:0] ? $signed(w_72) : $signed(_GEN_792); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_794 = 7'h49 == _temp_T_21[6:0] ? $signed(w_73) : $signed(_GEN_793); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_795 = 7'h4a == _temp_T_21[6:0] ? $signed(w_74) : $signed(_GEN_794); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_796 = 7'h4b == _temp_T_21[6:0] ? $signed(w_75) : $signed(_GEN_795); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_797 = 7'h4c == _temp_T_21[6:0] ? $signed(w_76) : $signed(_GEN_796); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_798 = 7'h4d == _temp_T_21[6:0] ? $signed(w_77) : $signed(_GEN_797); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_799 = 7'h4e == _temp_T_21[6:0] ? $signed(w_78) : $signed(_GEN_798); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_800 = 7'h4f == _temp_T_21[6:0] ? $signed(w_79) : $signed(_GEN_799); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_802 = 7'h1 == _temp_T_26[6:0] ? $signed(w_1) : $signed(w_0); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_803 = 7'h2 == _temp_T_26[6:0] ? $signed(w_2) : $signed(_GEN_802); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_804 = 7'h3 == _temp_T_26[6:0] ? $signed(w_3) : $signed(_GEN_803); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_805 = 7'h4 == _temp_T_26[6:0] ? $signed(w_4) : $signed(_GEN_804); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_806 = 7'h5 == _temp_T_26[6:0] ? $signed(w_5) : $signed(_GEN_805); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_807 = 7'h6 == _temp_T_26[6:0] ? $signed(w_6) : $signed(_GEN_806); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_808 = 7'h7 == _temp_T_26[6:0] ? $signed(w_7) : $signed(_GEN_807); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_809 = 7'h8 == _temp_T_26[6:0] ? $signed(w_8) : $signed(_GEN_808); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_810 = 7'h9 == _temp_T_26[6:0] ? $signed(w_9) : $signed(_GEN_809); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_811 = 7'ha == _temp_T_26[6:0] ? $signed(w_10) : $signed(_GEN_810); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_812 = 7'hb == _temp_T_26[6:0] ? $signed(w_11) : $signed(_GEN_811); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_813 = 7'hc == _temp_T_26[6:0] ? $signed(w_12) : $signed(_GEN_812); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_814 = 7'hd == _temp_T_26[6:0] ? $signed(w_13) : $signed(_GEN_813); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_815 = 7'he == _temp_T_26[6:0] ? $signed(w_14) : $signed(_GEN_814); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_816 = 7'hf == _temp_T_26[6:0] ? $signed(w_15) : $signed(_GEN_815); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_817 = 7'h10 == _temp_T_26[6:0] ? $signed(w_16) : $signed(_GEN_816); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_818 = 7'h11 == _temp_T_26[6:0] ? $signed(w_17) : $signed(_GEN_817); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_819 = 7'h12 == _temp_T_26[6:0] ? $signed(w_18) : $signed(_GEN_818); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_820 = 7'h13 == _temp_T_26[6:0] ? $signed(w_19) : $signed(_GEN_819); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_821 = 7'h14 == _temp_T_26[6:0] ? $signed(w_20) : $signed(_GEN_820); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_822 = 7'h15 == _temp_T_26[6:0] ? $signed(w_21) : $signed(_GEN_821); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_823 = 7'h16 == _temp_T_26[6:0] ? $signed(w_22) : $signed(_GEN_822); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_824 = 7'h17 == _temp_T_26[6:0] ? $signed(w_23) : $signed(_GEN_823); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_825 = 7'h18 == _temp_T_26[6:0] ? $signed(w_24) : $signed(_GEN_824); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_826 = 7'h19 == _temp_T_26[6:0] ? $signed(w_25) : $signed(_GEN_825); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_827 = 7'h1a == _temp_T_26[6:0] ? $signed(w_26) : $signed(_GEN_826); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_828 = 7'h1b == _temp_T_26[6:0] ? $signed(w_27) : $signed(_GEN_827); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_829 = 7'h1c == _temp_T_26[6:0] ? $signed(w_28) : $signed(_GEN_828); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_830 = 7'h1d == _temp_T_26[6:0] ? $signed(w_29) : $signed(_GEN_829); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_831 = 7'h1e == _temp_T_26[6:0] ? $signed(w_30) : $signed(_GEN_830); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_832 = 7'h1f == _temp_T_26[6:0] ? $signed(w_31) : $signed(_GEN_831); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_833 = 7'h20 == _temp_T_26[6:0] ? $signed(w_32) : $signed(_GEN_832); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_834 = 7'h21 == _temp_T_26[6:0] ? $signed(w_33) : $signed(_GEN_833); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_835 = 7'h22 == _temp_T_26[6:0] ? $signed(w_34) : $signed(_GEN_834); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_836 = 7'h23 == _temp_T_26[6:0] ? $signed(w_35) : $signed(_GEN_835); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_837 = 7'h24 == _temp_T_26[6:0] ? $signed(w_36) : $signed(_GEN_836); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_838 = 7'h25 == _temp_T_26[6:0] ? $signed(w_37) : $signed(_GEN_837); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_839 = 7'h26 == _temp_T_26[6:0] ? $signed(w_38) : $signed(_GEN_838); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_840 = 7'h27 == _temp_T_26[6:0] ? $signed(w_39) : $signed(_GEN_839); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_841 = 7'h28 == _temp_T_26[6:0] ? $signed(w_40) : $signed(_GEN_840); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_842 = 7'h29 == _temp_T_26[6:0] ? $signed(w_41) : $signed(_GEN_841); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_843 = 7'h2a == _temp_T_26[6:0] ? $signed(w_42) : $signed(_GEN_842); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_844 = 7'h2b == _temp_T_26[6:0] ? $signed(w_43) : $signed(_GEN_843); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_845 = 7'h2c == _temp_T_26[6:0] ? $signed(w_44) : $signed(_GEN_844); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_846 = 7'h2d == _temp_T_26[6:0] ? $signed(w_45) : $signed(_GEN_845); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_847 = 7'h2e == _temp_T_26[6:0] ? $signed(w_46) : $signed(_GEN_846); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_848 = 7'h2f == _temp_T_26[6:0] ? $signed(w_47) : $signed(_GEN_847); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_849 = 7'h30 == _temp_T_26[6:0] ? $signed(w_48) : $signed(_GEN_848); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_850 = 7'h31 == _temp_T_26[6:0] ? $signed(w_49) : $signed(_GEN_849); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_851 = 7'h32 == _temp_T_26[6:0] ? $signed(w_50) : $signed(_GEN_850); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_852 = 7'h33 == _temp_T_26[6:0] ? $signed(w_51) : $signed(_GEN_851); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_853 = 7'h34 == _temp_T_26[6:0] ? $signed(w_52) : $signed(_GEN_852); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_854 = 7'h35 == _temp_T_26[6:0] ? $signed(w_53) : $signed(_GEN_853); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_855 = 7'h36 == _temp_T_26[6:0] ? $signed(w_54) : $signed(_GEN_854); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_856 = 7'h37 == _temp_T_26[6:0] ? $signed(w_55) : $signed(_GEN_855); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_857 = 7'h38 == _temp_T_26[6:0] ? $signed(w_56) : $signed(_GEN_856); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_858 = 7'h39 == _temp_T_26[6:0] ? $signed(w_57) : $signed(_GEN_857); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_859 = 7'h3a == _temp_T_26[6:0] ? $signed(w_58) : $signed(_GEN_858); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_860 = 7'h3b == _temp_T_26[6:0] ? $signed(w_59) : $signed(_GEN_859); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_861 = 7'h3c == _temp_T_26[6:0] ? $signed(w_60) : $signed(_GEN_860); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_862 = 7'h3d == _temp_T_26[6:0] ? $signed(w_61) : $signed(_GEN_861); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_863 = 7'h3e == _temp_T_26[6:0] ? $signed(w_62) : $signed(_GEN_862); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_864 = 7'h3f == _temp_T_26[6:0] ? $signed(w_63) : $signed(_GEN_863); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_865 = 7'h40 == _temp_T_26[6:0] ? $signed(w_64) : $signed(_GEN_864); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_866 = 7'h41 == _temp_T_26[6:0] ? $signed(w_65) : $signed(_GEN_865); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_867 = 7'h42 == _temp_T_26[6:0] ? $signed(w_66) : $signed(_GEN_866); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_868 = 7'h43 == _temp_T_26[6:0] ? $signed(w_67) : $signed(_GEN_867); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_869 = 7'h44 == _temp_T_26[6:0] ? $signed(w_68) : $signed(_GEN_868); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_870 = 7'h45 == _temp_T_26[6:0] ? $signed(w_69) : $signed(_GEN_869); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_871 = 7'h46 == _temp_T_26[6:0] ? $signed(w_70) : $signed(_GEN_870); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_872 = 7'h47 == _temp_T_26[6:0] ? $signed(w_71) : $signed(_GEN_871); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_873 = 7'h48 == _temp_T_26[6:0] ? $signed(w_72) : $signed(_GEN_872); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_874 = 7'h49 == _temp_T_26[6:0] ? $signed(w_73) : $signed(_GEN_873); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_875 = 7'h4a == _temp_T_26[6:0] ? $signed(w_74) : $signed(_GEN_874); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_876 = 7'h4b == _temp_T_26[6:0] ? $signed(w_75) : $signed(_GEN_875); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_877 = 7'h4c == _temp_T_26[6:0] ? $signed(w_76) : $signed(_GEN_876); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_878 = 7'h4d == _temp_T_26[6:0] ? $signed(w_77) : $signed(_GEN_877); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_879 = 7'h4e == _temp_T_26[6:0] ? $signed(w_78) : $signed(_GEN_878); // @[digest.scala 186:{50,50}]
  wire [31:0] _GEN_880 = 7'h4f == _temp_T_26[6:0] ? $signed(w_79) : $signed(_GEN_879); // @[digest.scala 186:{50,50}]
  wire [31:0] _temp_T_29 = $signed(_GEN_800) ^ $signed(_GEN_880); // @[digest.scala 186:50]
  wire [31:0] _temp_T_33 = $signed(j) - 32'she; // @[digest.scala 186:109]
  wire [31:0] _GEN_882 = 7'h1 == _temp_T_33[6:0] ? $signed(w_1) : $signed(w_0); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_883 = 7'h2 == _temp_T_33[6:0] ? $signed(w_2) : $signed(_GEN_882); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_884 = 7'h3 == _temp_T_33[6:0] ? $signed(w_3) : $signed(_GEN_883); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_885 = 7'h4 == _temp_T_33[6:0] ? $signed(w_4) : $signed(_GEN_884); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_886 = 7'h5 == _temp_T_33[6:0] ? $signed(w_5) : $signed(_GEN_885); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_887 = 7'h6 == _temp_T_33[6:0] ? $signed(w_6) : $signed(_GEN_886); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_888 = 7'h7 == _temp_T_33[6:0] ? $signed(w_7) : $signed(_GEN_887); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_889 = 7'h8 == _temp_T_33[6:0] ? $signed(w_8) : $signed(_GEN_888); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_890 = 7'h9 == _temp_T_33[6:0] ? $signed(w_9) : $signed(_GEN_889); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_891 = 7'ha == _temp_T_33[6:0] ? $signed(w_10) : $signed(_GEN_890); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_892 = 7'hb == _temp_T_33[6:0] ? $signed(w_11) : $signed(_GEN_891); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_893 = 7'hc == _temp_T_33[6:0] ? $signed(w_12) : $signed(_GEN_892); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_894 = 7'hd == _temp_T_33[6:0] ? $signed(w_13) : $signed(_GEN_893); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_895 = 7'he == _temp_T_33[6:0] ? $signed(w_14) : $signed(_GEN_894); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_896 = 7'hf == _temp_T_33[6:0] ? $signed(w_15) : $signed(_GEN_895); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_897 = 7'h10 == _temp_T_33[6:0] ? $signed(w_16) : $signed(_GEN_896); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_898 = 7'h11 == _temp_T_33[6:0] ? $signed(w_17) : $signed(_GEN_897); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_899 = 7'h12 == _temp_T_33[6:0] ? $signed(w_18) : $signed(_GEN_898); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_900 = 7'h13 == _temp_T_33[6:0] ? $signed(w_19) : $signed(_GEN_899); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_901 = 7'h14 == _temp_T_33[6:0] ? $signed(w_20) : $signed(_GEN_900); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_902 = 7'h15 == _temp_T_33[6:0] ? $signed(w_21) : $signed(_GEN_901); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_903 = 7'h16 == _temp_T_33[6:0] ? $signed(w_22) : $signed(_GEN_902); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_904 = 7'h17 == _temp_T_33[6:0] ? $signed(w_23) : $signed(_GEN_903); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_905 = 7'h18 == _temp_T_33[6:0] ? $signed(w_24) : $signed(_GEN_904); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_906 = 7'h19 == _temp_T_33[6:0] ? $signed(w_25) : $signed(_GEN_905); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_907 = 7'h1a == _temp_T_33[6:0] ? $signed(w_26) : $signed(_GEN_906); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_908 = 7'h1b == _temp_T_33[6:0] ? $signed(w_27) : $signed(_GEN_907); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_909 = 7'h1c == _temp_T_33[6:0] ? $signed(w_28) : $signed(_GEN_908); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_910 = 7'h1d == _temp_T_33[6:0] ? $signed(w_29) : $signed(_GEN_909); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_911 = 7'h1e == _temp_T_33[6:0] ? $signed(w_30) : $signed(_GEN_910); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_912 = 7'h1f == _temp_T_33[6:0] ? $signed(w_31) : $signed(_GEN_911); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_913 = 7'h20 == _temp_T_33[6:0] ? $signed(w_32) : $signed(_GEN_912); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_914 = 7'h21 == _temp_T_33[6:0] ? $signed(w_33) : $signed(_GEN_913); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_915 = 7'h22 == _temp_T_33[6:0] ? $signed(w_34) : $signed(_GEN_914); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_916 = 7'h23 == _temp_T_33[6:0] ? $signed(w_35) : $signed(_GEN_915); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_917 = 7'h24 == _temp_T_33[6:0] ? $signed(w_36) : $signed(_GEN_916); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_918 = 7'h25 == _temp_T_33[6:0] ? $signed(w_37) : $signed(_GEN_917); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_919 = 7'h26 == _temp_T_33[6:0] ? $signed(w_38) : $signed(_GEN_918); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_920 = 7'h27 == _temp_T_33[6:0] ? $signed(w_39) : $signed(_GEN_919); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_921 = 7'h28 == _temp_T_33[6:0] ? $signed(w_40) : $signed(_GEN_920); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_922 = 7'h29 == _temp_T_33[6:0] ? $signed(w_41) : $signed(_GEN_921); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_923 = 7'h2a == _temp_T_33[6:0] ? $signed(w_42) : $signed(_GEN_922); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_924 = 7'h2b == _temp_T_33[6:0] ? $signed(w_43) : $signed(_GEN_923); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_925 = 7'h2c == _temp_T_33[6:0] ? $signed(w_44) : $signed(_GEN_924); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_926 = 7'h2d == _temp_T_33[6:0] ? $signed(w_45) : $signed(_GEN_925); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_927 = 7'h2e == _temp_T_33[6:0] ? $signed(w_46) : $signed(_GEN_926); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_928 = 7'h2f == _temp_T_33[6:0] ? $signed(w_47) : $signed(_GEN_927); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_929 = 7'h30 == _temp_T_33[6:0] ? $signed(w_48) : $signed(_GEN_928); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_930 = 7'h31 == _temp_T_33[6:0] ? $signed(w_49) : $signed(_GEN_929); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_931 = 7'h32 == _temp_T_33[6:0] ? $signed(w_50) : $signed(_GEN_930); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_932 = 7'h33 == _temp_T_33[6:0] ? $signed(w_51) : $signed(_GEN_931); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_933 = 7'h34 == _temp_T_33[6:0] ? $signed(w_52) : $signed(_GEN_932); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_934 = 7'h35 == _temp_T_33[6:0] ? $signed(w_53) : $signed(_GEN_933); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_935 = 7'h36 == _temp_T_33[6:0] ? $signed(w_54) : $signed(_GEN_934); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_936 = 7'h37 == _temp_T_33[6:0] ? $signed(w_55) : $signed(_GEN_935); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_937 = 7'h38 == _temp_T_33[6:0] ? $signed(w_56) : $signed(_GEN_936); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_938 = 7'h39 == _temp_T_33[6:0] ? $signed(w_57) : $signed(_GEN_937); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_939 = 7'h3a == _temp_T_33[6:0] ? $signed(w_58) : $signed(_GEN_938); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_940 = 7'h3b == _temp_T_33[6:0] ? $signed(w_59) : $signed(_GEN_939); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_941 = 7'h3c == _temp_T_33[6:0] ? $signed(w_60) : $signed(_GEN_940); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_942 = 7'h3d == _temp_T_33[6:0] ? $signed(w_61) : $signed(_GEN_941); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_943 = 7'h3e == _temp_T_33[6:0] ? $signed(w_62) : $signed(_GEN_942); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_944 = 7'h3f == _temp_T_33[6:0] ? $signed(w_63) : $signed(_GEN_943); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_945 = 7'h40 == _temp_T_33[6:0] ? $signed(w_64) : $signed(_GEN_944); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_946 = 7'h41 == _temp_T_33[6:0] ? $signed(w_65) : $signed(_GEN_945); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_947 = 7'h42 == _temp_T_33[6:0] ? $signed(w_66) : $signed(_GEN_946); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_948 = 7'h43 == _temp_T_33[6:0] ? $signed(w_67) : $signed(_GEN_947); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_949 = 7'h44 == _temp_T_33[6:0] ? $signed(w_68) : $signed(_GEN_948); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_950 = 7'h45 == _temp_T_33[6:0] ? $signed(w_69) : $signed(_GEN_949); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_951 = 7'h46 == _temp_T_33[6:0] ? $signed(w_70) : $signed(_GEN_950); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_952 = 7'h47 == _temp_T_33[6:0] ? $signed(w_71) : $signed(_GEN_951); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_953 = 7'h48 == _temp_T_33[6:0] ? $signed(w_72) : $signed(_GEN_952); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_954 = 7'h49 == _temp_T_33[6:0] ? $signed(w_73) : $signed(_GEN_953); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_955 = 7'h4a == _temp_T_33[6:0] ? $signed(w_74) : $signed(_GEN_954); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_956 = 7'h4b == _temp_T_33[6:0] ? $signed(w_75) : $signed(_GEN_955); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_957 = 7'h4c == _temp_T_33[6:0] ? $signed(w_76) : $signed(_GEN_956); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_958 = 7'h4d == _temp_T_33[6:0] ? $signed(w_77) : $signed(_GEN_957); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_959 = 7'h4e == _temp_T_33[6:0] ? $signed(w_78) : $signed(_GEN_958); // @[digest.scala 186:{81,81}]
  wire [31:0] _GEN_960 = 7'h4f == _temp_T_33[6:0] ? $signed(w_79) : $signed(_GEN_959); // @[digest.scala 186:{81,81}]
  wire [31:0] _temp_T_36 = $signed(_temp_T_29) ^ $signed(_GEN_960); // @[digest.scala 186:81]
  wire [31:0] _temp_T_40 = $signed(j) - 32'sh10; // @[digest.scala 186:141]
  wire [31:0] _GEN_962 = 7'h1 == _temp_T_40[6:0] ? $signed(w_1) : $signed(w_0); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_963 = 7'h2 == _temp_T_40[6:0] ? $signed(w_2) : $signed(_GEN_962); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_964 = 7'h3 == _temp_T_40[6:0] ? $signed(w_3) : $signed(_GEN_963); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_965 = 7'h4 == _temp_T_40[6:0] ? $signed(w_4) : $signed(_GEN_964); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_966 = 7'h5 == _temp_T_40[6:0] ? $signed(w_5) : $signed(_GEN_965); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_967 = 7'h6 == _temp_T_40[6:0] ? $signed(w_6) : $signed(_GEN_966); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_968 = 7'h7 == _temp_T_40[6:0] ? $signed(w_7) : $signed(_GEN_967); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_969 = 7'h8 == _temp_T_40[6:0] ? $signed(w_8) : $signed(_GEN_968); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_970 = 7'h9 == _temp_T_40[6:0] ? $signed(w_9) : $signed(_GEN_969); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_971 = 7'ha == _temp_T_40[6:0] ? $signed(w_10) : $signed(_GEN_970); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_972 = 7'hb == _temp_T_40[6:0] ? $signed(w_11) : $signed(_GEN_971); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_973 = 7'hc == _temp_T_40[6:0] ? $signed(w_12) : $signed(_GEN_972); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_974 = 7'hd == _temp_T_40[6:0] ? $signed(w_13) : $signed(_GEN_973); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_975 = 7'he == _temp_T_40[6:0] ? $signed(w_14) : $signed(_GEN_974); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_976 = 7'hf == _temp_T_40[6:0] ? $signed(w_15) : $signed(_GEN_975); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_977 = 7'h10 == _temp_T_40[6:0] ? $signed(w_16) : $signed(_GEN_976); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_978 = 7'h11 == _temp_T_40[6:0] ? $signed(w_17) : $signed(_GEN_977); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_979 = 7'h12 == _temp_T_40[6:0] ? $signed(w_18) : $signed(_GEN_978); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_980 = 7'h13 == _temp_T_40[6:0] ? $signed(w_19) : $signed(_GEN_979); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_981 = 7'h14 == _temp_T_40[6:0] ? $signed(w_20) : $signed(_GEN_980); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_982 = 7'h15 == _temp_T_40[6:0] ? $signed(w_21) : $signed(_GEN_981); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_983 = 7'h16 == _temp_T_40[6:0] ? $signed(w_22) : $signed(_GEN_982); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_984 = 7'h17 == _temp_T_40[6:0] ? $signed(w_23) : $signed(_GEN_983); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_985 = 7'h18 == _temp_T_40[6:0] ? $signed(w_24) : $signed(_GEN_984); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_986 = 7'h19 == _temp_T_40[6:0] ? $signed(w_25) : $signed(_GEN_985); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_987 = 7'h1a == _temp_T_40[6:0] ? $signed(w_26) : $signed(_GEN_986); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_988 = 7'h1b == _temp_T_40[6:0] ? $signed(w_27) : $signed(_GEN_987); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_989 = 7'h1c == _temp_T_40[6:0] ? $signed(w_28) : $signed(_GEN_988); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_990 = 7'h1d == _temp_T_40[6:0] ? $signed(w_29) : $signed(_GEN_989); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_991 = 7'h1e == _temp_T_40[6:0] ? $signed(w_30) : $signed(_GEN_990); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_992 = 7'h1f == _temp_T_40[6:0] ? $signed(w_31) : $signed(_GEN_991); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_993 = 7'h20 == _temp_T_40[6:0] ? $signed(w_32) : $signed(_GEN_992); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_994 = 7'h21 == _temp_T_40[6:0] ? $signed(w_33) : $signed(_GEN_993); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_995 = 7'h22 == _temp_T_40[6:0] ? $signed(w_34) : $signed(_GEN_994); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_996 = 7'h23 == _temp_T_40[6:0] ? $signed(w_35) : $signed(_GEN_995); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_997 = 7'h24 == _temp_T_40[6:0] ? $signed(w_36) : $signed(_GEN_996); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_998 = 7'h25 == _temp_T_40[6:0] ? $signed(w_37) : $signed(_GEN_997); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_999 = 7'h26 == _temp_T_40[6:0] ? $signed(w_38) : $signed(_GEN_998); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1000 = 7'h27 == _temp_T_40[6:0] ? $signed(w_39) : $signed(_GEN_999); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1001 = 7'h28 == _temp_T_40[6:0] ? $signed(w_40) : $signed(_GEN_1000); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1002 = 7'h29 == _temp_T_40[6:0] ? $signed(w_41) : $signed(_GEN_1001); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1003 = 7'h2a == _temp_T_40[6:0] ? $signed(w_42) : $signed(_GEN_1002); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1004 = 7'h2b == _temp_T_40[6:0] ? $signed(w_43) : $signed(_GEN_1003); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1005 = 7'h2c == _temp_T_40[6:0] ? $signed(w_44) : $signed(_GEN_1004); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1006 = 7'h2d == _temp_T_40[6:0] ? $signed(w_45) : $signed(_GEN_1005); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1007 = 7'h2e == _temp_T_40[6:0] ? $signed(w_46) : $signed(_GEN_1006); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1008 = 7'h2f == _temp_T_40[6:0] ? $signed(w_47) : $signed(_GEN_1007); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1009 = 7'h30 == _temp_T_40[6:0] ? $signed(w_48) : $signed(_GEN_1008); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1010 = 7'h31 == _temp_T_40[6:0] ? $signed(w_49) : $signed(_GEN_1009); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1011 = 7'h32 == _temp_T_40[6:0] ? $signed(w_50) : $signed(_GEN_1010); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1012 = 7'h33 == _temp_T_40[6:0] ? $signed(w_51) : $signed(_GEN_1011); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1013 = 7'h34 == _temp_T_40[6:0] ? $signed(w_52) : $signed(_GEN_1012); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1014 = 7'h35 == _temp_T_40[6:0] ? $signed(w_53) : $signed(_GEN_1013); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1015 = 7'h36 == _temp_T_40[6:0] ? $signed(w_54) : $signed(_GEN_1014); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1016 = 7'h37 == _temp_T_40[6:0] ? $signed(w_55) : $signed(_GEN_1015); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1017 = 7'h38 == _temp_T_40[6:0] ? $signed(w_56) : $signed(_GEN_1016); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1018 = 7'h39 == _temp_T_40[6:0] ? $signed(w_57) : $signed(_GEN_1017); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1019 = 7'h3a == _temp_T_40[6:0] ? $signed(w_58) : $signed(_GEN_1018); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1020 = 7'h3b == _temp_T_40[6:0] ? $signed(w_59) : $signed(_GEN_1019); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1021 = 7'h3c == _temp_T_40[6:0] ? $signed(w_60) : $signed(_GEN_1020); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1022 = 7'h3d == _temp_T_40[6:0] ? $signed(w_61) : $signed(_GEN_1021); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1023 = 7'h3e == _temp_T_40[6:0] ? $signed(w_62) : $signed(_GEN_1022); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1024 = 7'h3f == _temp_T_40[6:0] ? $signed(w_63) : $signed(_GEN_1023); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1025 = 7'h40 == _temp_T_40[6:0] ? $signed(w_64) : $signed(_GEN_1024); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1026 = 7'h41 == _temp_T_40[6:0] ? $signed(w_65) : $signed(_GEN_1025); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1027 = 7'h42 == _temp_T_40[6:0] ? $signed(w_66) : $signed(_GEN_1026); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1028 = 7'h43 == _temp_T_40[6:0] ? $signed(w_67) : $signed(_GEN_1027); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1029 = 7'h44 == _temp_T_40[6:0] ? $signed(w_68) : $signed(_GEN_1028); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1030 = 7'h45 == _temp_T_40[6:0] ? $signed(w_69) : $signed(_GEN_1029); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1031 = 7'h46 == _temp_T_40[6:0] ? $signed(w_70) : $signed(_GEN_1030); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1032 = 7'h47 == _temp_T_40[6:0] ? $signed(w_71) : $signed(_GEN_1031); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1033 = 7'h48 == _temp_T_40[6:0] ? $signed(w_72) : $signed(_GEN_1032); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1034 = 7'h49 == _temp_T_40[6:0] ? $signed(w_73) : $signed(_GEN_1033); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1035 = 7'h4a == _temp_T_40[6:0] ? $signed(w_74) : $signed(_GEN_1034); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1036 = 7'h4b == _temp_T_40[6:0] ? $signed(w_75) : $signed(_GEN_1035); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1037 = 7'h4c == _temp_T_40[6:0] ? $signed(w_76) : $signed(_GEN_1036); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1038 = 7'h4d == _temp_T_40[6:0] ? $signed(w_77) : $signed(_GEN_1037); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1039 = 7'h4e == _temp_T_40[6:0] ? $signed(w_78) : $signed(_GEN_1038); // @[digest.scala 186:{113,113}]
  wire [31:0] _GEN_1040 = 7'h4f == _temp_T_40[6:0] ? $signed(w_79) : $signed(_GEN_1039); // @[digest.scala 186:{113,113}]
  wire [31:0] _temp_T_43 = $signed(_temp_T_36) ^ $signed(_GEN_1040); // @[digest.scala 186:113]
  wire [31:0] _w_T_49 = __m_rol_0_io_out_rol; // @[digest.scala 190:{29,29}]
  wire [31:0] _GEN_1041 = 7'h0 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_0); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1042 = 7'h1 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_1); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1043 = 7'h2 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_2); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1044 = 7'h3 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_3); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1045 = 7'h4 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_4); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1046 = 7'h5 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_5); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1047 = 7'h6 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_6); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1048 = 7'h7 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_7); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1049 = 7'h8 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_8); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1050 = 7'h9 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_9); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1051 = 7'ha == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_10); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1052 = 7'hb == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_11); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1053 = 7'hc == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_12); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1054 = 7'hd == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_13); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1055 = 7'he == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_14); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1056 = 7'hf == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_15); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1057 = 7'h10 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_16); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1058 = 7'h11 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_17); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1059 = 7'h12 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_18); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1060 = 7'h13 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_19); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1061 = 7'h14 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_20); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1062 = 7'h15 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_21); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1063 = 7'h16 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_22); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1064 = 7'h17 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_23); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1065 = 7'h18 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_24); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1066 = 7'h19 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_25); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1067 = 7'h1a == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_26); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1068 = 7'h1b == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_27); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1069 = 7'h1c == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_28); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1070 = 7'h1d == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_29); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1071 = 7'h1e == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_30); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1072 = 7'h1f == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_31); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1073 = 7'h20 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_32); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1074 = 7'h21 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_33); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1075 = 7'h22 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_34); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1076 = 7'h23 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_35); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1077 = 7'h24 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_36); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1078 = 7'h25 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_37); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1079 = 7'h26 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_38); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1080 = 7'h27 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_39); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1081 = 7'h28 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_40); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1082 = 7'h29 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_41); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1083 = 7'h2a == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_42); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1084 = 7'h2b == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_43); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1085 = 7'h2c == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_44); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1086 = 7'h2d == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_45); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1087 = 7'h2e == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_46); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1088 = 7'h2f == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_47); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1089 = 7'h30 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_48); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1090 = 7'h31 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_49); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1091 = 7'h32 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_50); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1092 = 7'h33 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_51); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1093 = 7'h34 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_52); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1094 = 7'h35 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_53); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1095 = 7'h36 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_54); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1096 = 7'h37 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_55); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1097 = 7'h38 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_56); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1098 = 7'h39 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_57); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1099 = 7'h3a == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_58); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1100 = 7'h3b == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_59); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1101 = 7'h3c == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_60); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1102 = 7'h3d == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_61); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1103 = 7'h3e == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_62); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1104 = 7'h3f == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_63); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1105 = 7'h40 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_64); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1106 = 7'h41 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_65); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1107 = 7'h42 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_66); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1108 = 7'h43 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_67); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1109 = 7'h44 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_68); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1110 = 7'h45 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_69); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1111 = 7'h46 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_70); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1112 = 7'h47 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_71); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1113 = 7'h48 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_72); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1114 = 7'h49 == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_73); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1115 = 7'h4a == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_74); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1116 = 7'h4b == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_75); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1117 = 7'h4c == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_76); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1118 = 7'h4d == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_77); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1119 = 7'h4e == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_78); // @[digest.scala 190:{29,29} 40:16]
  wire [31:0] _GEN_1120 = 7'h4f == _T_44[6:0] ? $signed(_w_T_49) : $signed(w_79); // @[digest.scala 190:{29,29} 40:16]
  wire  __m_rol_0_io_valid_T = __m_rol_0_io_ready ? 1'h0 : 1'h1; // @[digest.scala 191:38]
  wire [5:0] _state_T_9 = __m_rol_0_io_ready ? 6'h1c : state; // @[digest.scala 194:25]
  wire [5:0] _state_T_11 = $signed(j) < 32'sh14 ? 6'h1d : 6'h20; // @[digest.scala 197:25]
  wire [31:0] _temp_T_45 = $signed(b) & $signed(c); // @[digest.scala 200:23]
  wire [31:0] _temp_T_47 = ~b; // @[digest.scala 204:29]
  wire [31:0] _temp_T_49 = $signed(_temp_T_47) & $signed(d); // @[digest.scala 204:33]
  wire [31:0] _temp_T_51 = $signed(temp) | $signed(_temp_T_49); // @[digest.scala 204:26]
  wire [31:0] _temp_T_54 = 32'sh5a827999 + $signed(temp); // @[digest.scala 208:41]
  wire [5:0] _state_T_13 = $signed(j) < 32'sh28 ? 6'h21 : 6'h23; // @[digest.scala 212:25]
  wire [31:0] _temp_T_56 = $signed(b) ^ $signed(c); // @[digest.scala 215:23]
  wire [31:0] _temp_T_58 = $signed(_temp_T_56) ^ $signed(d); // @[digest.scala 215:27]
  wire [31:0] _temp_T_61 = 32'sh6ed9eba1 + $signed(temp); // @[digest.scala 219:41]
  wire [5:0] _state_T_15 = $signed(j) < 32'sh3c ? 6'h24 : 6'h26; // @[digest.scala 223:25]
  wire [31:0] _temp_T_65 = $signed(b) & $signed(d); // @[digest.scala 226:31]
  wire [31:0] _temp_T_67 = $signed(_temp_T_45) | $signed(_temp_T_65); // @[digest.scala 226:27]
  wire [31:0] _temp_T_69 = $signed(c) & $signed(d); // @[digest.scala 226:39]
  wire [31:0] _temp_T_71 = $signed(_temp_T_67) | $signed(_temp_T_69); // @[digest.scala 226:35]
  wire [31:0] _temp_T_74 = $signed(temp) - 32'sh70e44324; // @[digest.scala 230:44]
  wire [31:0] _temp_T_81 = $signed(temp) - 32'sh359d3e2a; // @[digest.scala 238:43]
  wire  __m_rol_1_io_valid_T = __m_rol_1_io_ready ? 1'h0 : 1'h1; // @[digest.scala 243:38]
  wire [5:0] _state_T_16 = __m_rol_1_io_ready ? 6'h29 : state; // @[digest.scala 246:25]
  wire [31:0] _t_T_2 = $signed(t) + $signed(e); // @[digest.scala 249:20]
  wire [31:0] _GEN_1122 = 7'h1 == _T_44[6:0] ? $signed(w_1) : $signed(w_0); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1123 = 7'h2 == _T_44[6:0] ? $signed(w_2) : $signed(_GEN_1122); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1124 = 7'h3 == _T_44[6:0] ? $signed(w_3) : $signed(_GEN_1123); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1125 = 7'h4 == _T_44[6:0] ? $signed(w_4) : $signed(_GEN_1124); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1126 = 7'h5 == _T_44[6:0] ? $signed(w_5) : $signed(_GEN_1125); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1127 = 7'h6 == _T_44[6:0] ? $signed(w_6) : $signed(_GEN_1126); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1128 = 7'h7 == _T_44[6:0] ? $signed(w_7) : $signed(_GEN_1127); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1129 = 7'h8 == _T_44[6:0] ? $signed(w_8) : $signed(_GEN_1128); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1130 = 7'h9 == _T_44[6:0] ? $signed(w_9) : $signed(_GEN_1129); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1131 = 7'ha == _T_44[6:0] ? $signed(w_10) : $signed(_GEN_1130); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1132 = 7'hb == _T_44[6:0] ? $signed(w_11) : $signed(_GEN_1131); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1133 = 7'hc == _T_44[6:0] ? $signed(w_12) : $signed(_GEN_1132); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1134 = 7'hd == _T_44[6:0] ? $signed(w_13) : $signed(_GEN_1133); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1135 = 7'he == _T_44[6:0] ? $signed(w_14) : $signed(_GEN_1134); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1136 = 7'hf == _T_44[6:0] ? $signed(w_15) : $signed(_GEN_1135); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1137 = 7'h10 == _T_44[6:0] ? $signed(w_16) : $signed(_GEN_1136); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1138 = 7'h11 == _T_44[6:0] ? $signed(w_17) : $signed(_GEN_1137); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1139 = 7'h12 == _T_44[6:0] ? $signed(w_18) : $signed(_GEN_1138); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1140 = 7'h13 == _T_44[6:0] ? $signed(w_19) : $signed(_GEN_1139); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1141 = 7'h14 == _T_44[6:0] ? $signed(w_20) : $signed(_GEN_1140); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1142 = 7'h15 == _T_44[6:0] ? $signed(w_21) : $signed(_GEN_1141); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1143 = 7'h16 == _T_44[6:0] ? $signed(w_22) : $signed(_GEN_1142); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1144 = 7'h17 == _T_44[6:0] ? $signed(w_23) : $signed(_GEN_1143); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1145 = 7'h18 == _T_44[6:0] ? $signed(w_24) : $signed(_GEN_1144); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1146 = 7'h19 == _T_44[6:0] ? $signed(w_25) : $signed(_GEN_1145); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1147 = 7'h1a == _T_44[6:0] ? $signed(w_26) : $signed(_GEN_1146); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1148 = 7'h1b == _T_44[6:0] ? $signed(w_27) : $signed(_GEN_1147); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1149 = 7'h1c == _T_44[6:0] ? $signed(w_28) : $signed(_GEN_1148); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1150 = 7'h1d == _T_44[6:0] ? $signed(w_29) : $signed(_GEN_1149); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1151 = 7'h1e == _T_44[6:0] ? $signed(w_30) : $signed(_GEN_1150); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1152 = 7'h1f == _T_44[6:0] ? $signed(w_31) : $signed(_GEN_1151); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1153 = 7'h20 == _T_44[6:0] ? $signed(w_32) : $signed(_GEN_1152); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1154 = 7'h21 == _T_44[6:0] ? $signed(w_33) : $signed(_GEN_1153); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1155 = 7'h22 == _T_44[6:0] ? $signed(w_34) : $signed(_GEN_1154); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1156 = 7'h23 == _T_44[6:0] ? $signed(w_35) : $signed(_GEN_1155); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1157 = 7'h24 == _T_44[6:0] ? $signed(w_36) : $signed(_GEN_1156); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1158 = 7'h25 == _T_44[6:0] ? $signed(w_37) : $signed(_GEN_1157); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1159 = 7'h26 == _T_44[6:0] ? $signed(w_38) : $signed(_GEN_1158); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1160 = 7'h27 == _T_44[6:0] ? $signed(w_39) : $signed(_GEN_1159); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1161 = 7'h28 == _T_44[6:0] ? $signed(w_40) : $signed(_GEN_1160); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1162 = 7'h29 == _T_44[6:0] ? $signed(w_41) : $signed(_GEN_1161); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1163 = 7'h2a == _T_44[6:0] ? $signed(w_42) : $signed(_GEN_1162); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1164 = 7'h2b == _T_44[6:0] ? $signed(w_43) : $signed(_GEN_1163); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1165 = 7'h2c == _T_44[6:0] ? $signed(w_44) : $signed(_GEN_1164); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1166 = 7'h2d == _T_44[6:0] ? $signed(w_45) : $signed(_GEN_1165); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1167 = 7'h2e == _T_44[6:0] ? $signed(w_46) : $signed(_GEN_1166); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1168 = 7'h2f == _T_44[6:0] ? $signed(w_47) : $signed(_GEN_1167); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1169 = 7'h30 == _T_44[6:0] ? $signed(w_48) : $signed(_GEN_1168); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1170 = 7'h31 == _T_44[6:0] ? $signed(w_49) : $signed(_GEN_1169); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1171 = 7'h32 == _T_44[6:0] ? $signed(w_50) : $signed(_GEN_1170); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1172 = 7'h33 == _T_44[6:0] ? $signed(w_51) : $signed(_GEN_1171); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1173 = 7'h34 == _T_44[6:0] ? $signed(w_52) : $signed(_GEN_1172); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1174 = 7'h35 == _T_44[6:0] ? $signed(w_53) : $signed(_GEN_1173); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1175 = 7'h36 == _T_44[6:0] ? $signed(w_54) : $signed(_GEN_1174); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1176 = 7'h37 == _T_44[6:0] ? $signed(w_55) : $signed(_GEN_1175); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1177 = 7'h38 == _T_44[6:0] ? $signed(w_56) : $signed(_GEN_1176); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1178 = 7'h39 == _T_44[6:0] ? $signed(w_57) : $signed(_GEN_1177); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1179 = 7'h3a == _T_44[6:0] ? $signed(w_58) : $signed(_GEN_1178); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1180 = 7'h3b == _T_44[6:0] ? $signed(w_59) : $signed(_GEN_1179); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1181 = 7'h3c == _T_44[6:0] ? $signed(w_60) : $signed(_GEN_1180); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1182 = 7'h3d == _T_44[6:0] ? $signed(w_61) : $signed(_GEN_1181); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1183 = 7'h3e == _T_44[6:0] ? $signed(w_62) : $signed(_GEN_1182); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1184 = 7'h3f == _T_44[6:0] ? $signed(w_63) : $signed(_GEN_1183); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1185 = 7'h40 == _T_44[6:0] ? $signed(w_64) : $signed(_GEN_1184); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1186 = 7'h41 == _T_44[6:0] ? $signed(w_65) : $signed(_GEN_1185); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1187 = 7'h42 == _T_44[6:0] ? $signed(w_66) : $signed(_GEN_1186); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1188 = 7'h43 == _T_44[6:0] ? $signed(w_67) : $signed(_GEN_1187); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1189 = 7'h44 == _T_44[6:0] ? $signed(w_68) : $signed(_GEN_1188); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1190 = 7'h45 == _T_44[6:0] ? $signed(w_69) : $signed(_GEN_1189); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1191 = 7'h46 == _T_44[6:0] ? $signed(w_70) : $signed(_GEN_1190); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1192 = 7'h47 == _T_44[6:0] ? $signed(w_71) : $signed(_GEN_1191); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1193 = 7'h48 == _T_44[6:0] ? $signed(w_72) : $signed(_GEN_1192); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1194 = 7'h49 == _T_44[6:0] ? $signed(w_73) : $signed(_GEN_1193); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1195 = 7'h4a == _T_44[6:0] ? $signed(w_74) : $signed(_GEN_1194); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1196 = 7'h4b == _T_44[6:0] ? $signed(w_75) : $signed(_GEN_1195); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1197 = 7'h4c == _T_44[6:0] ? $signed(w_76) : $signed(_GEN_1196); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1198 = 7'h4d == _T_44[6:0] ? $signed(w_77) : $signed(_GEN_1197); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1199 = 7'h4e == _T_44[6:0] ? $signed(w_78) : $signed(_GEN_1198); // @[digest.scala 249:{24,24}]
  wire [31:0] _GEN_1200 = 7'h4f == _T_44[6:0] ? $signed(w_79) : $signed(_GEN_1199); // @[digest.scala 249:{24,24}]
  wire [31:0] _t_T_7 = $signed(_t_T_2) + $signed(_GEN_1200); // @[digest.scala 249:24]
  wire [31:0] _t_T_10 = $signed(_t_T_7) + $signed(temp); // @[digest.scala 249:42]
  wire  __m_rol_2_io_valid_T = __m_rol_2_io_ready ? 1'h0 : 1'h1; // @[digest.scala 262:38]
  wire [5:0] _state_T_17 = __m_rol_2_io_ready ? 6'h2d : state; // @[digest.scala 265:25]
  wire [31:0] _j_T_2 = $signed(j) + 32'sh1; // @[digest.scala 276:21]
  wire [31:0] _a_T_2 = $signed(a) + $signed(olda); // @[digest.scala 280:20]
  wire [31:0] _b_T_2 = $signed(b) + $signed(oldb); // @[digest.scala 284:20]
  wire [31:0] _c_T_2 = $signed(c) + $signed(oldc); // @[digest.scala 288:20]
  wire [31:0] _d_T_2 = $signed(d) + $signed(oldd); // @[digest.scala 292:20]
  wire [31:0] _e_T_2 = $signed(e) + $signed(olde); // @[digest.scala 296:20]
  wire [31:0] _i_T_5 = $signed(i) + 32'sh10; // @[digest.scala 300:20]
  wire [31:0] _GEN_1201 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_0) : $signed(digest_0); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1202 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_1) : $signed(digest_1); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1203 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_2) : $signed(digest_2); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1204 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_3) : $signed(digest_3); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1205 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_4) : $signed(digest_4); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1206 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_5) : $signed(digest_5); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1207 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_6) : $signed(digest_6); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1208 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_7) : $signed(digest_7); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1209 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_8) : $signed(digest_8); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1210 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_9) : $signed(digest_9); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1211 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_10) : $signed(digest_10); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1212 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_11) : $signed(digest_11); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1213 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_12) : $signed(digest_12); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1214 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_13) : $signed(digest_13); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1215 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_14) : $signed(digest_14); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1216 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_15) : $signed(digest_15); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1217 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_16) : $signed(digest_16); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1218 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_17) : $signed(digest_17); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1219 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_18) : $signed(digest_18); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1220 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_19) : $signed(digest_19); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1221 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_20) : $signed(digest_20); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1222 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_21) : $signed(digest_21); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1223 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_22) : $signed(digest_22); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1224 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_23) : $signed(digest_23); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1225 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_24) : $signed(digest_24); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1226 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_25) : $signed(digest_25); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1227 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_26) : $signed(digest_26); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1228 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_27) : $signed(digest_27); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1229 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_28) : $signed(digest_28); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1230 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_29) : $signed(digest_29); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1231 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_30) : $signed(digest_30); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1232 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_31) : $signed(digest_31); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1233 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_32) : $signed(digest_32); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1234 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_33) : $signed(digest_33); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1235 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_34) : $signed(digest_34); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1236 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_35) : $signed(digest_35); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1237 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_36) : $signed(digest_36); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1238 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_37) : $signed(digest_37); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1239 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_38) : $signed(digest_38); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1240 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_39) : $signed(digest_39); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1241 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_40) : $signed(digest_40); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1242 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_41) : $signed(digest_41); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1243 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_42) : $signed(digest_42); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1244 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_43) : $signed(digest_43); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1245 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_44) : $signed(digest_44); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1246 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_45) : $signed(digest_45); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1247 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_46) : $signed(digest_46); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1248 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_47) : $signed(digest_47); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1249 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_48) : $signed(digest_48); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1250 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_49) : $signed(digest_49); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1251 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_50) : $signed(digest_50); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1252 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_51) : $signed(digest_51); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1253 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_52) : $signed(digest_52); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1254 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_53) : $signed(digest_53); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1255 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_54) : $signed(digest_54); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1256 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_55) : $signed(digest_55); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1257 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_56) : $signed(digest_56); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1258 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_57) : $signed(digest_57); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1259 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_58) : $signed(digest_58); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1260 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_59) : $signed(digest_59); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1261 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_60) : $signed(digest_60); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1262 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_61) : $signed(digest_61); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1263 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_62) : $signed(digest_62); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1264 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_63) : $signed(digest_63); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1265 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_64) : $signed(digest_64); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1266 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_65) : $signed(digest_65); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1267 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_66) : $signed(digest_66); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1268 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_67) : $signed(digest_67); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1269 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_68) : $signed(digest_68); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1270 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_69) : $signed(digest_69); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1271 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_70) : $signed(digest_70); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1272 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_71) : $signed(digest_71); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1273 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_72) : $signed(digest_72); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1274 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_73) : $signed(digest_73); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1275 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_74) : $signed(digest_74); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1276 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_75) : $signed(digest_75); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1277 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_76) : $signed(digest_76); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1278 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_77) : $signed(digest_77); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1279 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_78) : $signed(digest_78); // @[digest.scala 306:38 307:24 53:21]
  wire [31:0] _GEN_1280 = __m_fill_0_io_ready ? $signed(__m_fill_0_io_arr_out_79) : $signed(digest_79); // @[digest.scala 306:38 307:24 53:21]
  wire  __m_fill_0_io_valid_T = __m_fill_0_io_ready ? 1'h0 : 1'h1; // @[digest.scala 310:39]
  wire [5:0] _state_T_18 = __m_fill_0_io_ready ? 6'h37 : state; // @[digest.scala 311:25]
  wire [31:0] _GEN_1281 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_0) : $signed(digest_0); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1282 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_1) : $signed(digest_1); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1283 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_2) : $signed(digest_2); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1284 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_3) : $signed(digest_3); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1285 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_4) : $signed(digest_4); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1286 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_5) : $signed(digest_5); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1287 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_6) : $signed(digest_6); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1288 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_7) : $signed(digest_7); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1289 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_8) : $signed(digest_8); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1290 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_9) : $signed(digest_9); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1291 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_10) : $signed(digest_10); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1292 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_11) : $signed(digest_11); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1293 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_12) : $signed(digest_12); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1294 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_13) : $signed(digest_13); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1295 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_14) : $signed(digest_14); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1296 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_15) : $signed(digest_15); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1297 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_16) : $signed(digest_16); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1298 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_17) : $signed(digest_17); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1299 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_18) : $signed(digest_18); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1300 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_19) : $signed(digest_19); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1301 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_20) : $signed(digest_20); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1302 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_21) : $signed(digest_21); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1303 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_22) : $signed(digest_22); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1304 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_23) : $signed(digest_23); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1305 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_24) : $signed(digest_24); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1306 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_25) : $signed(digest_25); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1307 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_26) : $signed(digest_26); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1308 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_27) : $signed(digest_27); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1309 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_28) : $signed(digest_28); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1310 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_29) : $signed(digest_29); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1311 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_30) : $signed(digest_30); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1312 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_31) : $signed(digest_31); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1313 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_32) : $signed(digest_32); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1314 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_33) : $signed(digest_33); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1315 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_34) : $signed(digest_34); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1316 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_35) : $signed(digest_35); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1317 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_36) : $signed(digest_36); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1318 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_37) : $signed(digest_37); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1319 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_38) : $signed(digest_38); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1320 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_39) : $signed(digest_39); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1321 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_40) : $signed(digest_40); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1322 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_41) : $signed(digest_41); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1323 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_42) : $signed(digest_42); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1324 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_43) : $signed(digest_43); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1325 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_44) : $signed(digest_44); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1326 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_45) : $signed(digest_45); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1327 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_46) : $signed(digest_46); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1328 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_47) : $signed(digest_47); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1329 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_48) : $signed(digest_48); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1330 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_49) : $signed(digest_49); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1331 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_50) : $signed(digest_50); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1332 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_51) : $signed(digest_51); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1333 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_52) : $signed(digest_52); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1334 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_53) : $signed(digest_53); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1335 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_54) : $signed(digest_54); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1336 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_55) : $signed(digest_55); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1337 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_56) : $signed(digest_56); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1338 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_57) : $signed(digest_57); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1339 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_58) : $signed(digest_58); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1340 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_59) : $signed(digest_59); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1341 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_60) : $signed(digest_60); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1342 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_61) : $signed(digest_61); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1343 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_62) : $signed(digest_62); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1344 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_63) : $signed(digest_63); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1345 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_64) : $signed(digest_64); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1346 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_65) : $signed(digest_65); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1347 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_66) : $signed(digest_66); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1348 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_67) : $signed(digest_67); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1349 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_68) : $signed(digest_68); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1350 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_69) : $signed(digest_69); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1351 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_70) : $signed(digest_70); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1352 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_71) : $signed(digest_71); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1353 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_72) : $signed(digest_72); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1354 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_73) : $signed(digest_73); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1355 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_74) : $signed(digest_74); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1356 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_75) : $signed(digest_75); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1357 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_76) : $signed(digest_76); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1358 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_77) : $signed(digest_77); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1359 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_78) : $signed(digest_78); // @[digest.scala 316:38 317:24 53:21]
  wire [31:0] _GEN_1360 = __m_fill_1_io_ready ? $signed(__m_fill_1_io_arr_out_79) : $signed(digest_79); // @[digest.scala 316:38 317:24 53:21]
  wire  __m_fill_1_io_valid_T = __m_fill_1_io_ready ? 1'h0 : 1'h1; // @[digest.scala 320:39]
  wire [5:0] _state_T_19 = __m_fill_1_io_ready ? 6'h38 : state; // @[digest.scala 321:25]
  wire [31:0] _GEN_1361 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_0) : $signed(digest_0); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1362 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_1) : $signed(digest_1); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1363 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_2) : $signed(digest_2); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1364 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_3) : $signed(digest_3); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1365 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_4) : $signed(digest_4); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1366 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_5) : $signed(digest_5); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1367 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_6) : $signed(digest_6); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1368 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_7) : $signed(digest_7); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1369 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_8) : $signed(digest_8); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1370 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_9) : $signed(digest_9); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1371 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_10) : $signed(digest_10); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1372 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_11) : $signed(digest_11); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1373 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_12) : $signed(digest_12); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1374 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_13) : $signed(digest_13); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1375 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_14) : $signed(digest_14); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1376 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_15) : $signed(digest_15); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1377 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_16) : $signed(digest_16); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1378 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_17) : $signed(digest_17); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1379 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_18) : $signed(digest_18); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1380 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_19) : $signed(digest_19); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1381 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_20) : $signed(digest_20); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1382 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_21) : $signed(digest_21); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1383 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_22) : $signed(digest_22); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1384 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_23) : $signed(digest_23); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1385 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_24) : $signed(digest_24); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1386 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_25) : $signed(digest_25); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1387 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_26) : $signed(digest_26); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1388 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_27) : $signed(digest_27); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1389 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_28) : $signed(digest_28); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1390 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_29) : $signed(digest_29); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1391 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_30) : $signed(digest_30); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1392 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_31) : $signed(digest_31); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1393 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_32) : $signed(digest_32); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1394 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_33) : $signed(digest_33); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1395 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_34) : $signed(digest_34); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1396 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_35) : $signed(digest_35); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1397 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_36) : $signed(digest_36); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1398 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_37) : $signed(digest_37); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1399 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_38) : $signed(digest_38); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1400 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_39) : $signed(digest_39); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1401 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_40) : $signed(digest_40); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1402 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_41) : $signed(digest_41); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1403 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_42) : $signed(digest_42); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1404 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_43) : $signed(digest_43); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1405 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_44) : $signed(digest_44); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1406 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_45) : $signed(digest_45); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1407 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_46) : $signed(digest_46); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1408 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_47) : $signed(digest_47); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1409 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_48) : $signed(digest_48); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1410 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_49) : $signed(digest_49); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1411 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_50) : $signed(digest_50); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1412 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_51) : $signed(digest_51); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1413 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_52) : $signed(digest_52); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1414 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_53) : $signed(digest_53); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1415 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_54) : $signed(digest_54); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1416 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_55) : $signed(digest_55); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1417 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_56) : $signed(digest_56); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1418 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_57) : $signed(digest_57); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1419 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_58) : $signed(digest_58); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1420 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_59) : $signed(digest_59); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1421 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_60) : $signed(digest_60); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1422 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_61) : $signed(digest_61); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1423 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_62) : $signed(digest_62); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1424 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_63) : $signed(digest_63); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1425 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_64) : $signed(digest_64); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1426 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_65) : $signed(digest_65); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1427 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_66) : $signed(digest_66); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1428 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_67) : $signed(digest_67); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1429 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_68) : $signed(digest_68); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1430 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_69) : $signed(digest_69); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1431 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_70) : $signed(digest_70); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1432 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_71) : $signed(digest_71); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1433 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_72) : $signed(digest_72); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1434 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_73) : $signed(digest_73); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1435 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_74) : $signed(digest_74); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1436 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_75) : $signed(digest_75); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1437 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_76) : $signed(digest_76); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1438 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_77) : $signed(digest_77); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1439 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_78) : $signed(digest_78); // @[digest.scala 326:38 327:24 53:21]
  wire [31:0] _GEN_1440 = __m_fill_2_io_ready ? $signed(__m_fill_2_io_arr_out_79) : $signed(digest_79); // @[digest.scala 326:38 327:24 53:21]
  wire  __m_fill_2_io_valid_T = __m_fill_2_io_ready ? 1'h0 : 1'h1; // @[digest.scala 330:39]
  wire [5:0] _state_T_20 = __m_fill_2_io_ready ? 6'h39 : state; // @[digest.scala 331:25]
  wire [31:0] _GEN_1441 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_0) : $signed(digest_0); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1442 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_1) : $signed(digest_1); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1443 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_2) : $signed(digest_2); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1444 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_3) : $signed(digest_3); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1445 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_4) : $signed(digest_4); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1446 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_5) : $signed(digest_5); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1447 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_6) : $signed(digest_6); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1448 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_7) : $signed(digest_7); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1449 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_8) : $signed(digest_8); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1450 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_9) : $signed(digest_9); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1451 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_10) : $signed(digest_10); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1452 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_11) : $signed(digest_11); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1453 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_12) : $signed(digest_12); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1454 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_13) : $signed(digest_13); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1455 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_14) : $signed(digest_14); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1456 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_15) : $signed(digest_15); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1457 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_16) : $signed(digest_16); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1458 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_17) : $signed(digest_17); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1459 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_18) : $signed(digest_18); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1460 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_19) : $signed(digest_19); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1461 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_20) : $signed(digest_20); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1462 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_21) : $signed(digest_21); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1463 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_22) : $signed(digest_22); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1464 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_23) : $signed(digest_23); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1465 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_24) : $signed(digest_24); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1466 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_25) : $signed(digest_25); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1467 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_26) : $signed(digest_26); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1468 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_27) : $signed(digest_27); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1469 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_28) : $signed(digest_28); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1470 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_29) : $signed(digest_29); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1471 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_30) : $signed(digest_30); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1472 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_31) : $signed(digest_31); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1473 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_32) : $signed(digest_32); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1474 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_33) : $signed(digest_33); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1475 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_34) : $signed(digest_34); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1476 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_35) : $signed(digest_35); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1477 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_36) : $signed(digest_36); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1478 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_37) : $signed(digest_37); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1479 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_38) : $signed(digest_38); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1480 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_39) : $signed(digest_39); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1481 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_40) : $signed(digest_40); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1482 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_41) : $signed(digest_41); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1483 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_42) : $signed(digest_42); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1484 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_43) : $signed(digest_43); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1485 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_44) : $signed(digest_44); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1486 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_45) : $signed(digest_45); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1487 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_46) : $signed(digest_46); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1488 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_47) : $signed(digest_47); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1489 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_48) : $signed(digest_48); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1490 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_49) : $signed(digest_49); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1491 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_50) : $signed(digest_50); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1492 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_51) : $signed(digest_51); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1493 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_52) : $signed(digest_52); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1494 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_53) : $signed(digest_53); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1495 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_54) : $signed(digest_54); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1496 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_55) : $signed(digest_55); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1497 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_56) : $signed(digest_56); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1498 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_57) : $signed(digest_57); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1499 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_58) : $signed(digest_58); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1500 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_59) : $signed(digest_59); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1501 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_60) : $signed(digest_60); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1502 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_61) : $signed(digest_61); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1503 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_62) : $signed(digest_62); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1504 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_63) : $signed(digest_63); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1505 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_64) : $signed(digest_64); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1506 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_65) : $signed(digest_65); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1507 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_66) : $signed(digest_66); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1508 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_67) : $signed(digest_67); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1509 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_68) : $signed(digest_68); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1510 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_69) : $signed(digest_69); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1511 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_70) : $signed(digest_70); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1512 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_71) : $signed(digest_71); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1513 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_72) : $signed(digest_72); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1514 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_73) : $signed(digest_73); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1515 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_74) : $signed(digest_74); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1516 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_75) : $signed(digest_75); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1517 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_76) : $signed(digest_76); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1518 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_77) : $signed(digest_77); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1519 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_78) : $signed(digest_78); // @[digest.scala 336:38 337:24 53:21]
  wire [31:0] _GEN_1520 = __m_fill_3_io_ready ? $signed(__m_fill_3_io_arr_out_79) : $signed(digest_79); // @[digest.scala 336:38 337:24 53:21]
  wire  __m_fill_3_io_valid_T = __m_fill_3_io_ready ? 1'h0 : 1'h1; // @[digest.scala 340:39]
  wire [5:0] _state_T_21 = __m_fill_3_io_ready ? 6'h3a : state; // @[digest.scala 341:25]
  wire [31:0] _GEN_1521 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_0) : $signed(digest_0); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1522 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_1) : $signed(digest_1); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1523 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_2) : $signed(digest_2); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1524 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_3) : $signed(digest_3); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1525 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_4) : $signed(digest_4); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1526 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_5) : $signed(digest_5); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1527 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_6) : $signed(digest_6); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1528 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_7) : $signed(digest_7); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1529 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_8) : $signed(digest_8); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1530 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_9) : $signed(digest_9); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1531 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_10) : $signed(digest_10); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1532 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_11) : $signed(digest_11); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1533 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_12) : $signed(digest_12); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1534 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_13) : $signed(digest_13); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1535 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_14) : $signed(digest_14); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1536 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_15) : $signed(digest_15); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1537 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_16) : $signed(digest_16); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1538 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_17) : $signed(digest_17); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1539 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_18) : $signed(digest_18); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1540 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_19) : $signed(digest_19); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1541 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_20) : $signed(digest_20); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1542 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_21) : $signed(digest_21); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1543 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_22) : $signed(digest_22); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1544 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_23) : $signed(digest_23); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1545 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_24) : $signed(digest_24); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1546 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_25) : $signed(digest_25); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1547 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_26) : $signed(digest_26); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1548 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_27) : $signed(digest_27); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1549 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_28) : $signed(digest_28); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1550 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_29) : $signed(digest_29); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1551 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_30) : $signed(digest_30); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1552 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_31) : $signed(digest_31); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1553 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_32) : $signed(digest_32); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1554 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_33) : $signed(digest_33); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1555 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_34) : $signed(digest_34); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1556 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_35) : $signed(digest_35); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1557 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_36) : $signed(digest_36); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1558 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_37) : $signed(digest_37); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1559 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_38) : $signed(digest_38); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1560 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_39) : $signed(digest_39); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1561 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_40) : $signed(digest_40); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1562 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_41) : $signed(digest_41); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1563 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_42) : $signed(digest_42); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1564 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_43) : $signed(digest_43); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1565 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_44) : $signed(digest_44); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1566 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_45) : $signed(digest_45); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1567 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_46) : $signed(digest_46); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1568 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_47) : $signed(digest_47); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1569 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_48) : $signed(digest_48); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1570 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_49) : $signed(digest_49); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1571 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_50) : $signed(digest_50); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1572 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_51) : $signed(digest_51); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1573 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_52) : $signed(digest_52); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1574 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_53) : $signed(digest_53); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1575 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_54) : $signed(digest_54); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1576 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_55) : $signed(digest_55); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1577 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_56) : $signed(digest_56); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1578 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_57) : $signed(digest_57); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1579 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_58) : $signed(digest_58); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1580 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_59) : $signed(digest_59); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1581 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_60) : $signed(digest_60); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1582 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_61) : $signed(digest_61); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1583 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_62) : $signed(digest_62); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1584 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_63) : $signed(digest_63); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1585 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_64) : $signed(digest_64); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1586 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_65) : $signed(digest_65); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1587 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_66) : $signed(digest_66); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1588 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_67) : $signed(digest_67); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1589 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_68) : $signed(digest_68); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1590 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_69) : $signed(digest_69); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1591 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_70) : $signed(digest_70); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1592 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_71) : $signed(digest_71); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1593 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_72) : $signed(digest_72); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1594 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_73) : $signed(digest_73); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1595 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_74) : $signed(digest_74); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1596 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_75) : $signed(digest_75); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1597 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_76) : $signed(digest_76); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1598 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_77) : $signed(digest_77); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1599 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_78) : $signed(digest_78); // @[digest.scala 346:38 347:24 53:21]
  wire [31:0] _GEN_1600 = __m_fill_4_io_ready ? $signed(__m_fill_4_io_arr_out_79) : $signed(digest_79); // @[digest.scala 346:38 347:24 53:21]
  wire  __m_fill_4_io_valid_T = __m_fill_4_io_ready ? 1'h0 : 1'h1; // @[digest.scala 350:39]
  wire [5:0] _state_T_22 = __m_fill_4_io_ready ? 6'h3b : state; // @[digest.scala 351:25]
  wire [5:0] _GEN_1601 = 6'h3b == state ? 6'h3f : _GEN_0; // @[digest.scala 354:19 81:19]
  wire [31:0] _GEN_1683 = 6'h3a == state ? $signed(_GEN_1521) : $signed(digest_0); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1684 = 6'h3a == state ? $signed(_GEN_1522) : $signed(digest_1); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1685 = 6'h3a == state ? $signed(_GEN_1523) : $signed(digest_2); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1686 = 6'h3a == state ? $signed(_GEN_1524) : $signed(digest_3); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1687 = 6'h3a == state ? $signed(_GEN_1525) : $signed(digest_4); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1688 = 6'h3a == state ? $signed(_GEN_1526) : $signed(digest_5); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1689 = 6'h3a == state ? $signed(_GEN_1527) : $signed(digest_6); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1690 = 6'h3a == state ? $signed(_GEN_1528) : $signed(digest_7); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1691 = 6'h3a == state ? $signed(_GEN_1529) : $signed(digest_8); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1692 = 6'h3a == state ? $signed(_GEN_1530) : $signed(digest_9); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1693 = 6'h3a == state ? $signed(_GEN_1531) : $signed(digest_10); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1694 = 6'h3a == state ? $signed(_GEN_1532) : $signed(digest_11); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1695 = 6'h3a == state ? $signed(_GEN_1533) : $signed(digest_12); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1696 = 6'h3a == state ? $signed(_GEN_1534) : $signed(digest_13); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1697 = 6'h3a == state ? $signed(_GEN_1535) : $signed(digest_14); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1698 = 6'h3a == state ? $signed(_GEN_1536) : $signed(digest_15); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1699 = 6'h3a == state ? $signed(_GEN_1537) : $signed(digest_16); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1700 = 6'h3a == state ? $signed(_GEN_1538) : $signed(digest_17); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1701 = 6'h3a == state ? $signed(_GEN_1539) : $signed(digest_18); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1702 = 6'h3a == state ? $signed(_GEN_1540) : $signed(digest_19); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1703 = 6'h3a == state ? $signed(_GEN_1541) : $signed(digest_20); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1704 = 6'h3a == state ? $signed(_GEN_1542) : $signed(digest_21); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1705 = 6'h3a == state ? $signed(_GEN_1543) : $signed(digest_22); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1706 = 6'h3a == state ? $signed(_GEN_1544) : $signed(digest_23); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1707 = 6'h3a == state ? $signed(_GEN_1545) : $signed(digest_24); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1708 = 6'h3a == state ? $signed(_GEN_1546) : $signed(digest_25); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1709 = 6'h3a == state ? $signed(_GEN_1547) : $signed(digest_26); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1710 = 6'h3a == state ? $signed(_GEN_1548) : $signed(digest_27); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1711 = 6'h3a == state ? $signed(_GEN_1549) : $signed(digest_28); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1712 = 6'h3a == state ? $signed(_GEN_1550) : $signed(digest_29); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1713 = 6'h3a == state ? $signed(_GEN_1551) : $signed(digest_30); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1714 = 6'h3a == state ? $signed(_GEN_1552) : $signed(digest_31); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1715 = 6'h3a == state ? $signed(_GEN_1553) : $signed(digest_32); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1716 = 6'h3a == state ? $signed(_GEN_1554) : $signed(digest_33); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1717 = 6'h3a == state ? $signed(_GEN_1555) : $signed(digest_34); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1718 = 6'h3a == state ? $signed(_GEN_1556) : $signed(digest_35); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1719 = 6'h3a == state ? $signed(_GEN_1557) : $signed(digest_36); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1720 = 6'h3a == state ? $signed(_GEN_1558) : $signed(digest_37); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1721 = 6'h3a == state ? $signed(_GEN_1559) : $signed(digest_38); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1722 = 6'h3a == state ? $signed(_GEN_1560) : $signed(digest_39); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1723 = 6'h3a == state ? $signed(_GEN_1561) : $signed(digest_40); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1724 = 6'h3a == state ? $signed(_GEN_1562) : $signed(digest_41); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1725 = 6'h3a == state ? $signed(_GEN_1563) : $signed(digest_42); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1726 = 6'h3a == state ? $signed(_GEN_1564) : $signed(digest_43); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1727 = 6'h3a == state ? $signed(_GEN_1565) : $signed(digest_44); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1728 = 6'h3a == state ? $signed(_GEN_1566) : $signed(digest_45); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1729 = 6'h3a == state ? $signed(_GEN_1567) : $signed(digest_46); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1730 = 6'h3a == state ? $signed(_GEN_1568) : $signed(digest_47); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1731 = 6'h3a == state ? $signed(_GEN_1569) : $signed(digest_48); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1732 = 6'h3a == state ? $signed(_GEN_1570) : $signed(digest_49); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1733 = 6'h3a == state ? $signed(_GEN_1571) : $signed(digest_50); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1734 = 6'h3a == state ? $signed(_GEN_1572) : $signed(digest_51); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1735 = 6'h3a == state ? $signed(_GEN_1573) : $signed(digest_52); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1736 = 6'h3a == state ? $signed(_GEN_1574) : $signed(digest_53); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1737 = 6'h3a == state ? $signed(_GEN_1575) : $signed(digest_54); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1738 = 6'h3a == state ? $signed(_GEN_1576) : $signed(digest_55); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1739 = 6'h3a == state ? $signed(_GEN_1577) : $signed(digest_56); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1740 = 6'h3a == state ? $signed(_GEN_1578) : $signed(digest_57); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1741 = 6'h3a == state ? $signed(_GEN_1579) : $signed(digest_58); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1742 = 6'h3a == state ? $signed(_GEN_1580) : $signed(digest_59); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1743 = 6'h3a == state ? $signed(_GEN_1581) : $signed(digest_60); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1744 = 6'h3a == state ? $signed(_GEN_1582) : $signed(digest_61); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1745 = 6'h3a == state ? $signed(_GEN_1583) : $signed(digest_62); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1746 = 6'h3a == state ? $signed(_GEN_1584) : $signed(digest_63); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1747 = 6'h3a == state ? $signed(_GEN_1585) : $signed(digest_64); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1748 = 6'h3a == state ? $signed(_GEN_1586) : $signed(digest_65); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1749 = 6'h3a == state ? $signed(_GEN_1587) : $signed(digest_66); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1750 = 6'h3a == state ? $signed(_GEN_1588) : $signed(digest_67); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1751 = 6'h3a == state ? $signed(_GEN_1589) : $signed(digest_68); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1752 = 6'h3a == state ? $signed(_GEN_1590) : $signed(digest_69); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1753 = 6'h3a == state ? $signed(_GEN_1591) : $signed(digest_70); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1754 = 6'h3a == state ? $signed(_GEN_1592) : $signed(digest_71); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1755 = 6'h3a == state ? $signed(_GEN_1593) : $signed(digest_72); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1756 = 6'h3a == state ? $signed(_GEN_1594) : $signed(digest_73); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1757 = 6'h3a == state ? $signed(_GEN_1595) : $signed(digest_74); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1758 = 6'h3a == state ? $signed(_GEN_1596) : $signed(digest_75); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1759 = 6'h3a == state ? $signed(_GEN_1597) : $signed(digest_76); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1760 = 6'h3a == state ? $signed(_GEN_1598) : $signed(digest_77); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1761 = 6'h3a == state ? $signed(_GEN_1599) : $signed(digest_78); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_1762 = 6'h3a == state ? $signed(_GEN_1600) : $signed(digest_79); // @[digest.scala 81:19 53:21]
  wire  _GEN_1764 = 6'h3a == state & __m_fill_4_io_valid_T; // @[digest.scala 81:19 350:33 78:25]
  wire [5:0] _GEN_1765 = 6'h3a == state ? _state_T_22 : _GEN_1601; // @[digest.scala 351:19 81:19]
  wire [31:0] _GEN_1847 = 6'h39 == state ? $signed(_GEN_1441) : $signed(_GEN_1683); // @[digest.scala 81:19]
  wire [31:0] _GEN_1848 = 6'h39 == state ? $signed(_GEN_1442) : $signed(_GEN_1684); // @[digest.scala 81:19]
  wire [31:0] _GEN_1849 = 6'h39 == state ? $signed(_GEN_1443) : $signed(_GEN_1685); // @[digest.scala 81:19]
  wire [31:0] _GEN_1850 = 6'h39 == state ? $signed(_GEN_1444) : $signed(_GEN_1686); // @[digest.scala 81:19]
  wire [31:0] _GEN_1851 = 6'h39 == state ? $signed(_GEN_1445) : $signed(_GEN_1687); // @[digest.scala 81:19]
  wire [31:0] _GEN_1852 = 6'h39 == state ? $signed(_GEN_1446) : $signed(_GEN_1688); // @[digest.scala 81:19]
  wire [31:0] _GEN_1853 = 6'h39 == state ? $signed(_GEN_1447) : $signed(_GEN_1689); // @[digest.scala 81:19]
  wire [31:0] _GEN_1854 = 6'h39 == state ? $signed(_GEN_1448) : $signed(_GEN_1690); // @[digest.scala 81:19]
  wire [31:0] _GEN_1855 = 6'h39 == state ? $signed(_GEN_1449) : $signed(_GEN_1691); // @[digest.scala 81:19]
  wire [31:0] _GEN_1856 = 6'h39 == state ? $signed(_GEN_1450) : $signed(_GEN_1692); // @[digest.scala 81:19]
  wire [31:0] _GEN_1857 = 6'h39 == state ? $signed(_GEN_1451) : $signed(_GEN_1693); // @[digest.scala 81:19]
  wire [31:0] _GEN_1858 = 6'h39 == state ? $signed(_GEN_1452) : $signed(_GEN_1694); // @[digest.scala 81:19]
  wire [31:0] _GEN_1859 = 6'h39 == state ? $signed(_GEN_1453) : $signed(_GEN_1695); // @[digest.scala 81:19]
  wire [31:0] _GEN_1860 = 6'h39 == state ? $signed(_GEN_1454) : $signed(_GEN_1696); // @[digest.scala 81:19]
  wire [31:0] _GEN_1861 = 6'h39 == state ? $signed(_GEN_1455) : $signed(_GEN_1697); // @[digest.scala 81:19]
  wire [31:0] _GEN_1862 = 6'h39 == state ? $signed(_GEN_1456) : $signed(_GEN_1698); // @[digest.scala 81:19]
  wire [31:0] _GEN_1863 = 6'h39 == state ? $signed(_GEN_1457) : $signed(_GEN_1699); // @[digest.scala 81:19]
  wire [31:0] _GEN_1864 = 6'h39 == state ? $signed(_GEN_1458) : $signed(_GEN_1700); // @[digest.scala 81:19]
  wire [31:0] _GEN_1865 = 6'h39 == state ? $signed(_GEN_1459) : $signed(_GEN_1701); // @[digest.scala 81:19]
  wire [31:0] _GEN_1866 = 6'h39 == state ? $signed(_GEN_1460) : $signed(_GEN_1702); // @[digest.scala 81:19]
  wire [31:0] _GEN_1867 = 6'h39 == state ? $signed(_GEN_1461) : $signed(_GEN_1703); // @[digest.scala 81:19]
  wire [31:0] _GEN_1868 = 6'h39 == state ? $signed(_GEN_1462) : $signed(_GEN_1704); // @[digest.scala 81:19]
  wire [31:0] _GEN_1869 = 6'h39 == state ? $signed(_GEN_1463) : $signed(_GEN_1705); // @[digest.scala 81:19]
  wire [31:0] _GEN_1870 = 6'h39 == state ? $signed(_GEN_1464) : $signed(_GEN_1706); // @[digest.scala 81:19]
  wire [31:0] _GEN_1871 = 6'h39 == state ? $signed(_GEN_1465) : $signed(_GEN_1707); // @[digest.scala 81:19]
  wire [31:0] _GEN_1872 = 6'h39 == state ? $signed(_GEN_1466) : $signed(_GEN_1708); // @[digest.scala 81:19]
  wire [31:0] _GEN_1873 = 6'h39 == state ? $signed(_GEN_1467) : $signed(_GEN_1709); // @[digest.scala 81:19]
  wire [31:0] _GEN_1874 = 6'h39 == state ? $signed(_GEN_1468) : $signed(_GEN_1710); // @[digest.scala 81:19]
  wire [31:0] _GEN_1875 = 6'h39 == state ? $signed(_GEN_1469) : $signed(_GEN_1711); // @[digest.scala 81:19]
  wire [31:0] _GEN_1876 = 6'h39 == state ? $signed(_GEN_1470) : $signed(_GEN_1712); // @[digest.scala 81:19]
  wire [31:0] _GEN_1877 = 6'h39 == state ? $signed(_GEN_1471) : $signed(_GEN_1713); // @[digest.scala 81:19]
  wire [31:0] _GEN_1878 = 6'h39 == state ? $signed(_GEN_1472) : $signed(_GEN_1714); // @[digest.scala 81:19]
  wire [31:0] _GEN_1879 = 6'h39 == state ? $signed(_GEN_1473) : $signed(_GEN_1715); // @[digest.scala 81:19]
  wire [31:0] _GEN_1880 = 6'h39 == state ? $signed(_GEN_1474) : $signed(_GEN_1716); // @[digest.scala 81:19]
  wire [31:0] _GEN_1881 = 6'h39 == state ? $signed(_GEN_1475) : $signed(_GEN_1717); // @[digest.scala 81:19]
  wire [31:0] _GEN_1882 = 6'h39 == state ? $signed(_GEN_1476) : $signed(_GEN_1718); // @[digest.scala 81:19]
  wire [31:0] _GEN_1883 = 6'h39 == state ? $signed(_GEN_1477) : $signed(_GEN_1719); // @[digest.scala 81:19]
  wire [31:0] _GEN_1884 = 6'h39 == state ? $signed(_GEN_1478) : $signed(_GEN_1720); // @[digest.scala 81:19]
  wire [31:0] _GEN_1885 = 6'h39 == state ? $signed(_GEN_1479) : $signed(_GEN_1721); // @[digest.scala 81:19]
  wire [31:0] _GEN_1886 = 6'h39 == state ? $signed(_GEN_1480) : $signed(_GEN_1722); // @[digest.scala 81:19]
  wire [31:0] _GEN_1887 = 6'h39 == state ? $signed(_GEN_1481) : $signed(_GEN_1723); // @[digest.scala 81:19]
  wire [31:0] _GEN_1888 = 6'h39 == state ? $signed(_GEN_1482) : $signed(_GEN_1724); // @[digest.scala 81:19]
  wire [31:0] _GEN_1889 = 6'h39 == state ? $signed(_GEN_1483) : $signed(_GEN_1725); // @[digest.scala 81:19]
  wire [31:0] _GEN_1890 = 6'h39 == state ? $signed(_GEN_1484) : $signed(_GEN_1726); // @[digest.scala 81:19]
  wire [31:0] _GEN_1891 = 6'h39 == state ? $signed(_GEN_1485) : $signed(_GEN_1727); // @[digest.scala 81:19]
  wire [31:0] _GEN_1892 = 6'h39 == state ? $signed(_GEN_1486) : $signed(_GEN_1728); // @[digest.scala 81:19]
  wire [31:0] _GEN_1893 = 6'h39 == state ? $signed(_GEN_1487) : $signed(_GEN_1729); // @[digest.scala 81:19]
  wire [31:0] _GEN_1894 = 6'h39 == state ? $signed(_GEN_1488) : $signed(_GEN_1730); // @[digest.scala 81:19]
  wire [31:0] _GEN_1895 = 6'h39 == state ? $signed(_GEN_1489) : $signed(_GEN_1731); // @[digest.scala 81:19]
  wire [31:0] _GEN_1896 = 6'h39 == state ? $signed(_GEN_1490) : $signed(_GEN_1732); // @[digest.scala 81:19]
  wire [31:0] _GEN_1897 = 6'h39 == state ? $signed(_GEN_1491) : $signed(_GEN_1733); // @[digest.scala 81:19]
  wire [31:0] _GEN_1898 = 6'h39 == state ? $signed(_GEN_1492) : $signed(_GEN_1734); // @[digest.scala 81:19]
  wire [31:0] _GEN_1899 = 6'h39 == state ? $signed(_GEN_1493) : $signed(_GEN_1735); // @[digest.scala 81:19]
  wire [31:0] _GEN_1900 = 6'h39 == state ? $signed(_GEN_1494) : $signed(_GEN_1736); // @[digest.scala 81:19]
  wire [31:0] _GEN_1901 = 6'h39 == state ? $signed(_GEN_1495) : $signed(_GEN_1737); // @[digest.scala 81:19]
  wire [31:0] _GEN_1902 = 6'h39 == state ? $signed(_GEN_1496) : $signed(_GEN_1738); // @[digest.scala 81:19]
  wire [31:0] _GEN_1903 = 6'h39 == state ? $signed(_GEN_1497) : $signed(_GEN_1739); // @[digest.scala 81:19]
  wire [31:0] _GEN_1904 = 6'h39 == state ? $signed(_GEN_1498) : $signed(_GEN_1740); // @[digest.scala 81:19]
  wire [31:0] _GEN_1905 = 6'h39 == state ? $signed(_GEN_1499) : $signed(_GEN_1741); // @[digest.scala 81:19]
  wire [31:0] _GEN_1906 = 6'h39 == state ? $signed(_GEN_1500) : $signed(_GEN_1742); // @[digest.scala 81:19]
  wire [31:0] _GEN_1907 = 6'h39 == state ? $signed(_GEN_1501) : $signed(_GEN_1743); // @[digest.scala 81:19]
  wire [31:0] _GEN_1908 = 6'h39 == state ? $signed(_GEN_1502) : $signed(_GEN_1744); // @[digest.scala 81:19]
  wire [31:0] _GEN_1909 = 6'h39 == state ? $signed(_GEN_1503) : $signed(_GEN_1745); // @[digest.scala 81:19]
  wire [31:0] _GEN_1910 = 6'h39 == state ? $signed(_GEN_1504) : $signed(_GEN_1746); // @[digest.scala 81:19]
  wire [31:0] _GEN_1911 = 6'h39 == state ? $signed(_GEN_1505) : $signed(_GEN_1747); // @[digest.scala 81:19]
  wire [31:0] _GEN_1912 = 6'h39 == state ? $signed(_GEN_1506) : $signed(_GEN_1748); // @[digest.scala 81:19]
  wire [31:0] _GEN_1913 = 6'h39 == state ? $signed(_GEN_1507) : $signed(_GEN_1749); // @[digest.scala 81:19]
  wire [31:0] _GEN_1914 = 6'h39 == state ? $signed(_GEN_1508) : $signed(_GEN_1750); // @[digest.scala 81:19]
  wire [31:0] _GEN_1915 = 6'h39 == state ? $signed(_GEN_1509) : $signed(_GEN_1751); // @[digest.scala 81:19]
  wire [31:0] _GEN_1916 = 6'h39 == state ? $signed(_GEN_1510) : $signed(_GEN_1752); // @[digest.scala 81:19]
  wire [31:0] _GEN_1917 = 6'h39 == state ? $signed(_GEN_1511) : $signed(_GEN_1753); // @[digest.scala 81:19]
  wire [31:0] _GEN_1918 = 6'h39 == state ? $signed(_GEN_1512) : $signed(_GEN_1754); // @[digest.scala 81:19]
  wire [31:0] _GEN_1919 = 6'h39 == state ? $signed(_GEN_1513) : $signed(_GEN_1755); // @[digest.scala 81:19]
  wire [31:0] _GEN_1920 = 6'h39 == state ? $signed(_GEN_1514) : $signed(_GEN_1756); // @[digest.scala 81:19]
  wire [31:0] _GEN_1921 = 6'h39 == state ? $signed(_GEN_1515) : $signed(_GEN_1757); // @[digest.scala 81:19]
  wire [31:0] _GEN_1922 = 6'h39 == state ? $signed(_GEN_1516) : $signed(_GEN_1758); // @[digest.scala 81:19]
  wire [31:0] _GEN_1923 = 6'h39 == state ? $signed(_GEN_1517) : $signed(_GEN_1759); // @[digest.scala 81:19]
  wire [31:0] _GEN_1924 = 6'h39 == state ? $signed(_GEN_1518) : $signed(_GEN_1760); // @[digest.scala 81:19]
  wire [31:0] _GEN_1925 = 6'h39 == state ? $signed(_GEN_1519) : $signed(_GEN_1761); // @[digest.scala 81:19]
  wire [31:0] _GEN_1926 = 6'h39 == state ? $signed(_GEN_1520) : $signed(_GEN_1762); // @[digest.scala 81:19]
  wire  _GEN_1928 = 6'h39 == state & __m_fill_3_io_valid_T; // @[digest.scala 81:19 340:33 73:25]
  wire [5:0] _GEN_1929 = 6'h39 == state ? _state_T_21 : _GEN_1765; // @[digest.scala 341:19 81:19]
  wire  _GEN_2012 = 6'h39 == state ? 1'h0 : _GEN_1764; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_2094 = 6'h38 == state ? $signed(_GEN_1361) : $signed(_GEN_1847); // @[digest.scala 81:19]
  wire [31:0] _GEN_2095 = 6'h38 == state ? $signed(_GEN_1362) : $signed(_GEN_1848); // @[digest.scala 81:19]
  wire [31:0] _GEN_2096 = 6'h38 == state ? $signed(_GEN_1363) : $signed(_GEN_1849); // @[digest.scala 81:19]
  wire [31:0] _GEN_2097 = 6'h38 == state ? $signed(_GEN_1364) : $signed(_GEN_1850); // @[digest.scala 81:19]
  wire [31:0] _GEN_2098 = 6'h38 == state ? $signed(_GEN_1365) : $signed(_GEN_1851); // @[digest.scala 81:19]
  wire [31:0] _GEN_2099 = 6'h38 == state ? $signed(_GEN_1366) : $signed(_GEN_1852); // @[digest.scala 81:19]
  wire [31:0] _GEN_2100 = 6'h38 == state ? $signed(_GEN_1367) : $signed(_GEN_1853); // @[digest.scala 81:19]
  wire [31:0] _GEN_2101 = 6'h38 == state ? $signed(_GEN_1368) : $signed(_GEN_1854); // @[digest.scala 81:19]
  wire [31:0] _GEN_2102 = 6'h38 == state ? $signed(_GEN_1369) : $signed(_GEN_1855); // @[digest.scala 81:19]
  wire [31:0] _GEN_2103 = 6'h38 == state ? $signed(_GEN_1370) : $signed(_GEN_1856); // @[digest.scala 81:19]
  wire [31:0] _GEN_2104 = 6'h38 == state ? $signed(_GEN_1371) : $signed(_GEN_1857); // @[digest.scala 81:19]
  wire [31:0] _GEN_2105 = 6'h38 == state ? $signed(_GEN_1372) : $signed(_GEN_1858); // @[digest.scala 81:19]
  wire [31:0] _GEN_2106 = 6'h38 == state ? $signed(_GEN_1373) : $signed(_GEN_1859); // @[digest.scala 81:19]
  wire [31:0] _GEN_2107 = 6'h38 == state ? $signed(_GEN_1374) : $signed(_GEN_1860); // @[digest.scala 81:19]
  wire [31:0] _GEN_2108 = 6'h38 == state ? $signed(_GEN_1375) : $signed(_GEN_1861); // @[digest.scala 81:19]
  wire [31:0] _GEN_2109 = 6'h38 == state ? $signed(_GEN_1376) : $signed(_GEN_1862); // @[digest.scala 81:19]
  wire [31:0] _GEN_2110 = 6'h38 == state ? $signed(_GEN_1377) : $signed(_GEN_1863); // @[digest.scala 81:19]
  wire [31:0] _GEN_2111 = 6'h38 == state ? $signed(_GEN_1378) : $signed(_GEN_1864); // @[digest.scala 81:19]
  wire [31:0] _GEN_2112 = 6'h38 == state ? $signed(_GEN_1379) : $signed(_GEN_1865); // @[digest.scala 81:19]
  wire [31:0] _GEN_2113 = 6'h38 == state ? $signed(_GEN_1380) : $signed(_GEN_1866); // @[digest.scala 81:19]
  wire [31:0] _GEN_2114 = 6'h38 == state ? $signed(_GEN_1381) : $signed(_GEN_1867); // @[digest.scala 81:19]
  wire [31:0] _GEN_2115 = 6'h38 == state ? $signed(_GEN_1382) : $signed(_GEN_1868); // @[digest.scala 81:19]
  wire [31:0] _GEN_2116 = 6'h38 == state ? $signed(_GEN_1383) : $signed(_GEN_1869); // @[digest.scala 81:19]
  wire [31:0] _GEN_2117 = 6'h38 == state ? $signed(_GEN_1384) : $signed(_GEN_1870); // @[digest.scala 81:19]
  wire [31:0] _GEN_2118 = 6'h38 == state ? $signed(_GEN_1385) : $signed(_GEN_1871); // @[digest.scala 81:19]
  wire [31:0] _GEN_2119 = 6'h38 == state ? $signed(_GEN_1386) : $signed(_GEN_1872); // @[digest.scala 81:19]
  wire [31:0] _GEN_2120 = 6'h38 == state ? $signed(_GEN_1387) : $signed(_GEN_1873); // @[digest.scala 81:19]
  wire [31:0] _GEN_2121 = 6'h38 == state ? $signed(_GEN_1388) : $signed(_GEN_1874); // @[digest.scala 81:19]
  wire [31:0] _GEN_2122 = 6'h38 == state ? $signed(_GEN_1389) : $signed(_GEN_1875); // @[digest.scala 81:19]
  wire [31:0] _GEN_2123 = 6'h38 == state ? $signed(_GEN_1390) : $signed(_GEN_1876); // @[digest.scala 81:19]
  wire [31:0] _GEN_2124 = 6'h38 == state ? $signed(_GEN_1391) : $signed(_GEN_1877); // @[digest.scala 81:19]
  wire [31:0] _GEN_2125 = 6'h38 == state ? $signed(_GEN_1392) : $signed(_GEN_1878); // @[digest.scala 81:19]
  wire [31:0] _GEN_2126 = 6'h38 == state ? $signed(_GEN_1393) : $signed(_GEN_1879); // @[digest.scala 81:19]
  wire [31:0] _GEN_2127 = 6'h38 == state ? $signed(_GEN_1394) : $signed(_GEN_1880); // @[digest.scala 81:19]
  wire [31:0] _GEN_2128 = 6'h38 == state ? $signed(_GEN_1395) : $signed(_GEN_1881); // @[digest.scala 81:19]
  wire [31:0] _GEN_2129 = 6'h38 == state ? $signed(_GEN_1396) : $signed(_GEN_1882); // @[digest.scala 81:19]
  wire [31:0] _GEN_2130 = 6'h38 == state ? $signed(_GEN_1397) : $signed(_GEN_1883); // @[digest.scala 81:19]
  wire [31:0] _GEN_2131 = 6'h38 == state ? $signed(_GEN_1398) : $signed(_GEN_1884); // @[digest.scala 81:19]
  wire [31:0] _GEN_2132 = 6'h38 == state ? $signed(_GEN_1399) : $signed(_GEN_1885); // @[digest.scala 81:19]
  wire [31:0] _GEN_2133 = 6'h38 == state ? $signed(_GEN_1400) : $signed(_GEN_1886); // @[digest.scala 81:19]
  wire [31:0] _GEN_2134 = 6'h38 == state ? $signed(_GEN_1401) : $signed(_GEN_1887); // @[digest.scala 81:19]
  wire [31:0] _GEN_2135 = 6'h38 == state ? $signed(_GEN_1402) : $signed(_GEN_1888); // @[digest.scala 81:19]
  wire [31:0] _GEN_2136 = 6'h38 == state ? $signed(_GEN_1403) : $signed(_GEN_1889); // @[digest.scala 81:19]
  wire [31:0] _GEN_2137 = 6'h38 == state ? $signed(_GEN_1404) : $signed(_GEN_1890); // @[digest.scala 81:19]
  wire [31:0] _GEN_2138 = 6'h38 == state ? $signed(_GEN_1405) : $signed(_GEN_1891); // @[digest.scala 81:19]
  wire [31:0] _GEN_2139 = 6'h38 == state ? $signed(_GEN_1406) : $signed(_GEN_1892); // @[digest.scala 81:19]
  wire [31:0] _GEN_2140 = 6'h38 == state ? $signed(_GEN_1407) : $signed(_GEN_1893); // @[digest.scala 81:19]
  wire [31:0] _GEN_2141 = 6'h38 == state ? $signed(_GEN_1408) : $signed(_GEN_1894); // @[digest.scala 81:19]
  wire [31:0] _GEN_2142 = 6'h38 == state ? $signed(_GEN_1409) : $signed(_GEN_1895); // @[digest.scala 81:19]
  wire [31:0] _GEN_2143 = 6'h38 == state ? $signed(_GEN_1410) : $signed(_GEN_1896); // @[digest.scala 81:19]
  wire [31:0] _GEN_2144 = 6'h38 == state ? $signed(_GEN_1411) : $signed(_GEN_1897); // @[digest.scala 81:19]
  wire [31:0] _GEN_2145 = 6'h38 == state ? $signed(_GEN_1412) : $signed(_GEN_1898); // @[digest.scala 81:19]
  wire [31:0] _GEN_2146 = 6'h38 == state ? $signed(_GEN_1413) : $signed(_GEN_1899); // @[digest.scala 81:19]
  wire [31:0] _GEN_2147 = 6'h38 == state ? $signed(_GEN_1414) : $signed(_GEN_1900); // @[digest.scala 81:19]
  wire [31:0] _GEN_2148 = 6'h38 == state ? $signed(_GEN_1415) : $signed(_GEN_1901); // @[digest.scala 81:19]
  wire [31:0] _GEN_2149 = 6'h38 == state ? $signed(_GEN_1416) : $signed(_GEN_1902); // @[digest.scala 81:19]
  wire [31:0] _GEN_2150 = 6'h38 == state ? $signed(_GEN_1417) : $signed(_GEN_1903); // @[digest.scala 81:19]
  wire [31:0] _GEN_2151 = 6'h38 == state ? $signed(_GEN_1418) : $signed(_GEN_1904); // @[digest.scala 81:19]
  wire [31:0] _GEN_2152 = 6'h38 == state ? $signed(_GEN_1419) : $signed(_GEN_1905); // @[digest.scala 81:19]
  wire [31:0] _GEN_2153 = 6'h38 == state ? $signed(_GEN_1420) : $signed(_GEN_1906); // @[digest.scala 81:19]
  wire [31:0] _GEN_2154 = 6'h38 == state ? $signed(_GEN_1421) : $signed(_GEN_1907); // @[digest.scala 81:19]
  wire [31:0] _GEN_2155 = 6'h38 == state ? $signed(_GEN_1422) : $signed(_GEN_1908); // @[digest.scala 81:19]
  wire [31:0] _GEN_2156 = 6'h38 == state ? $signed(_GEN_1423) : $signed(_GEN_1909); // @[digest.scala 81:19]
  wire [31:0] _GEN_2157 = 6'h38 == state ? $signed(_GEN_1424) : $signed(_GEN_1910); // @[digest.scala 81:19]
  wire [31:0] _GEN_2158 = 6'h38 == state ? $signed(_GEN_1425) : $signed(_GEN_1911); // @[digest.scala 81:19]
  wire [31:0] _GEN_2159 = 6'h38 == state ? $signed(_GEN_1426) : $signed(_GEN_1912); // @[digest.scala 81:19]
  wire [31:0] _GEN_2160 = 6'h38 == state ? $signed(_GEN_1427) : $signed(_GEN_1913); // @[digest.scala 81:19]
  wire [31:0] _GEN_2161 = 6'h38 == state ? $signed(_GEN_1428) : $signed(_GEN_1914); // @[digest.scala 81:19]
  wire [31:0] _GEN_2162 = 6'h38 == state ? $signed(_GEN_1429) : $signed(_GEN_1915); // @[digest.scala 81:19]
  wire [31:0] _GEN_2163 = 6'h38 == state ? $signed(_GEN_1430) : $signed(_GEN_1916); // @[digest.scala 81:19]
  wire [31:0] _GEN_2164 = 6'h38 == state ? $signed(_GEN_1431) : $signed(_GEN_1917); // @[digest.scala 81:19]
  wire [31:0] _GEN_2165 = 6'h38 == state ? $signed(_GEN_1432) : $signed(_GEN_1918); // @[digest.scala 81:19]
  wire [31:0] _GEN_2166 = 6'h38 == state ? $signed(_GEN_1433) : $signed(_GEN_1919); // @[digest.scala 81:19]
  wire [31:0] _GEN_2167 = 6'h38 == state ? $signed(_GEN_1434) : $signed(_GEN_1920); // @[digest.scala 81:19]
  wire [31:0] _GEN_2168 = 6'h38 == state ? $signed(_GEN_1435) : $signed(_GEN_1921); // @[digest.scala 81:19]
  wire [31:0] _GEN_2169 = 6'h38 == state ? $signed(_GEN_1436) : $signed(_GEN_1922); // @[digest.scala 81:19]
  wire [31:0] _GEN_2170 = 6'h38 == state ? $signed(_GEN_1437) : $signed(_GEN_1923); // @[digest.scala 81:19]
  wire [31:0] _GEN_2171 = 6'h38 == state ? $signed(_GEN_1438) : $signed(_GEN_1924); // @[digest.scala 81:19]
  wire [31:0] _GEN_2172 = 6'h38 == state ? $signed(_GEN_1439) : $signed(_GEN_1925); // @[digest.scala 81:19]
  wire [31:0] _GEN_2173 = 6'h38 == state ? $signed(_GEN_1440) : $signed(_GEN_1926); // @[digest.scala 81:19]
  wire  _GEN_2175 = 6'h38 == state & __m_fill_2_io_valid_T; // @[digest.scala 81:19 330:33 68:25]
  wire [5:0] _GEN_2176 = 6'h38 == state ? _state_T_20 : _GEN_1929; // @[digest.scala 331:19 81:19]
  wire  _GEN_2259 = 6'h38 == state ? 1'h0 : _GEN_1928; // @[digest.scala 81:19 73:25]
  wire  _GEN_2342 = 6'h38 == state ? 1'h0 : _GEN_2012; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_2424 = 6'h37 == state ? $signed(_GEN_1281) : $signed(_GEN_2094); // @[digest.scala 81:19]
  wire [31:0] _GEN_2425 = 6'h37 == state ? $signed(_GEN_1282) : $signed(_GEN_2095); // @[digest.scala 81:19]
  wire [31:0] _GEN_2426 = 6'h37 == state ? $signed(_GEN_1283) : $signed(_GEN_2096); // @[digest.scala 81:19]
  wire [31:0] _GEN_2427 = 6'h37 == state ? $signed(_GEN_1284) : $signed(_GEN_2097); // @[digest.scala 81:19]
  wire [31:0] _GEN_2428 = 6'h37 == state ? $signed(_GEN_1285) : $signed(_GEN_2098); // @[digest.scala 81:19]
  wire [31:0] _GEN_2429 = 6'h37 == state ? $signed(_GEN_1286) : $signed(_GEN_2099); // @[digest.scala 81:19]
  wire [31:0] _GEN_2430 = 6'h37 == state ? $signed(_GEN_1287) : $signed(_GEN_2100); // @[digest.scala 81:19]
  wire [31:0] _GEN_2431 = 6'h37 == state ? $signed(_GEN_1288) : $signed(_GEN_2101); // @[digest.scala 81:19]
  wire [31:0] _GEN_2432 = 6'h37 == state ? $signed(_GEN_1289) : $signed(_GEN_2102); // @[digest.scala 81:19]
  wire [31:0] _GEN_2433 = 6'h37 == state ? $signed(_GEN_1290) : $signed(_GEN_2103); // @[digest.scala 81:19]
  wire [31:0] _GEN_2434 = 6'h37 == state ? $signed(_GEN_1291) : $signed(_GEN_2104); // @[digest.scala 81:19]
  wire [31:0] _GEN_2435 = 6'h37 == state ? $signed(_GEN_1292) : $signed(_GEN_2105); // @[digest.scala 81:19]
  wire [31:0] _GEN_2436 = 6'h37 == state ? $signed(_GEN_1293) : $signed(_GEN_2106); // @[digest.scala 81:19]
  wire [31:0] _GEN_2437 = 6'h37 == state ? $signed(_GEN_1294) : $signed(_GEN_2107); // @[digest.scala 81:19]
  wire [31:0] _GEN_2438 = 6'h37 == state ? $signed(_GEN_1295) : $signed(_GEN_2108); // @[digest.scala 81:19]
  wire [31:0] _GEN_2439 = 6'h37 == state ? $signed(_GEN_1296) : $signed(_GEN_2109); // @[digest.scala 81:19]
  wire [31:0] _GEN_2440 = 6'h37 == state ? $signed(_GEN_1297) : $signed(_GEN_2110); // @[digest.scala 81:19]
  wire [31:0] _GEN_2441 = 6'h37 == state ? $signed(_GEN_1298) : $signed(_GEN_2111); // @[digest.scala 81:19]
  wire [31:0] _GEN_2442 = 6'h37 == state ? $signed(_GEN_1299) : $signed(_GEN_2112); // @[digest.scala 81:19]
  wire [31:0] _GEN_2443 = 6'h37 == state ? $signed(_GEN_1300) : $signed(_GEN_2113); // @[digest.scala 81:19]
  wire [31:0] _GEN_2444 = 6'h37 == state ? $signed(_GEN_1301) : $signed(_GEN_2114); // @[digest.scala 81:19]
  wire [31:0] _GEN_2445 = 6'h37 == state ? $signed(_GEN_1302) : $signed(_GEN_2115); // @[digest.scala 81:19]
  wire [31:0] _GEN_2446 = 6'h37 == state ? $signed(_GEN_1303) : $signed(_GEN_2116); // @[digest.scala 81:19]
  wire [31:0] _GEN_2447 = 6'h37 == state ? $signed(_GEN_1304) : $signed(_GEN_2117); // @[digest.scala 81:19]
  wire [31:0] _GEN_2448 = 6'h37 == state ? $signed(_GEN_1305) : $signed(_GEN_2118); // @[digest.scala 81:19]
  wire [31:0] _GEN_2449 = 6'h37 == state ? $signed(_GEN_1306) : $signed(_GEN_2119); // @[digest.scala 81:19]
  wire [31:0] _GEN_2450 = 6'h37 == state ? $signed(_GEN_1307) : $signed(_GEN_2120); // @[digest.scala 81:19]
  wire [31:0] _GEN_2451 = 6'h37 == state ? $signed(_GEN_1308) : $signed(_GEN_2121); // @[digest.scala 81:19]
  wire [31:0] _GEN_2452 = 6'h37 == state ? $signed(_GEN_1309) : $signed(_GEN_2122); // @[digest.scala 81:19]
  wire [31:0] _GEN_2453 = 6'h37 == state ? $signed(_GEN_1310) : $signed(_GEN_2123); // @[digest.scala 81:19]
  wire [31:0] _GEN_2454 = 6'h37 == state ? $signed(_GEN_1311) : $signed(_GEN_2124); // @[digest.scala 81:19]
  wire [31:0] _GEN_2455 = 6'h37 == state ? $signed(_GEN_1312) : $signed(_GEN_2125); // @[digest.scala 81:19]
  wire [31:0] _GEN_2456 = 6'h37 == state ? $signed(_GEN_1313) : $signed(_GEN_2126); // @[digest.scala 81:19]
  wire [31:0] _GEN_2457 = 6'h37 == state ? $signed(_GEN_1314) : $signed(_GEN_2127); // @[digest.scala 81:19]
  wire [31:0] _GEN_2458 = 6'h37 == state ? $signed(_GEN_1315) : $signed(_GEN_2128); // @[digest.scala 81:19]
  wire [31:0] _GEN_2459 = 6'h37 == state ? $signed(_GEN_1316) : $signed(_GEN_2129); // @[digest.scala 81:19]
  wire [31:0] _GEN_2460 = 6'h37 == state ? $signed(_GEN_1317) : $signed(_GEN_2130); // @[digest.scala 81:19]
  wire [31:0] _GEN_2461 = 6'h37 == state ? $signed(_GEN_1318) : $signed(_GEN_2131); // @[digest.scala 81:19]
  wire [31:0] _GEN_2462 = 6'h37 == state ? $signed(_GEN_1319) : $signed(_GEN_2132); // @[digest.scala 81:19]
  wire [31:0] _GEN_2463 = 6'h37 == state ? $signed(_GEN_1320) : $signed(_GEN_2133); // @[digest.scala 81:19]
  wire [31:0] _GEN_2464 = 6'h37 == state ? $signed(_GEN_1321) : $signed(_GEN_2134); // @[digest.scala 81:19]
  wire [31:0] _GEN_2465 = 6'h37 == state ? $signed(_GEN_1322) : $signed(_GEN_2135); // @[digest.scala 81:19]
  wire [31:0] _GEN_2466 = 6'h37 == state ? $signed(_GEN_1323) : $signed(_GEN_2136); // @[digest.scala 81:19]
  wire [31:0] _GEN_2467 = 6'h37 == state ? $signed(_GEN_1324) : $signed(_GEN_2137); // @[digest.scala 81:19]
  wire [31:0] _GEN_2468 = 6'h37 == state ? $signed(_GEN_1325) : $signed(_GEN_2138); // @[digest.scala 81:19]
  wire [31:0] _GEN_2469 = 6'h37 == state ? $signed(_GEN_1326) : $signed(_GEN_2139); // @[digest.scala 81:19]
  wire [31:0] _GEN_2470 = 6'h37 == state ? $signed(_GEN_1327) : $signed(_GEN_2140); // @[digest.scala 81:19]
  wire [31:0] _GEN_2471 = 6'h37 == state ? $signed(_GEN_1328) : $signed(_GEN_2141); // @[digest.scala 81:19]
  wire [31:0] _GEN_2472 = 6'h37 == state ? $signed(_GEN_1329) : $signed(_GEN_2142); // @[digest.scala 81:19]
  wire [31:0] _GEN_2473 = 6'h37 == state ? $signed(_GEN_1330) : $signed(_GEN_2143); // @[digest.scala 81:19]
  wire [31:0] _GEN_2474 = 6'h37 == state ? $signed(_GEN_1331) : $signed(_GEN_2144); // @[digest.scala 81:19]
  wire [31:0] _GEN_2475 = 6'h37 == state ? $signed(_GEN_1332) : $signed(_GEN_2145); // @[digest.scala 81:19]
  wire [31:0] _GEN_2476 = 6'h37 == state ? $signed(_GEN_1333) : $signed(_GEN_2146); // @[digest.scala 81:19]
  wire [31:0] _GEN_2477 = 6'h37 == state ? $signed(_GEN_1334) : $signed(_GEN_2147); // @[digest.scala 81:19]
  wire [31:0] _GEN_2478 = 6'h37 == state ? $signed(_GEN_1335) : $signed(_GEN_2148); // @[digest.scala 81:19]
  wire [31:0] _GEN_2479 = 6'h37 == state ? $signed(_GEN_1336) : $signed(_GEN_2149); // @[digest.scala 81:19]
  wire [31:0] _GEN_2480 = 6'h37 == state ? $signed(_GEN_1337) : $signed(_GEN_2150); // @[digest.scala 81:19]
  wire [31:0] _GEN_2481 = 6'h37 == state ? $signed(_GEN_1338) : $signed(_GEN_2151); // @[digest.scala 81:19]
  wire [31:0] _GEN_2482 = 6'h37 == state ? $signed(_GEN_1339) : $signed(_GEN_2152); // @[digest.scala 81:19]
  wire [31:0] _GEN_2483 = 6'h37 == state ? $signed(_GEN_1340) : $signed(_GEN_2153); // @[digest.scala 81:19]
  wire [31:0] _GEN_2484 = 6'h37 == state ? $signed(_GEN_1341) : $signed(_GEN_2154); // @[digest.scala 81:19]
  wire [31:0] _GEN_2485 = 6'h37 == state ? $signed(_GEN_1342) : $signed(_GEN_2155); // @[digest.scala 81:19]
  wire [31:0] _GEN_2486 = 6'h37 == state ? $signed(_GEN_1343) : $signed(_GEN_2156); // @[digest.scala 81:19]
  wire [31:0] _GEN_2487 = 6'h37 == state ? $signed(_GEN_1344) : $signed(_GEN_2157); // @[digest.scala 81:19]
  wire [31:0] _GEN_2488 = 6'h37 == state ? $signed(_GEN_1345) : $signed(_GEN_2158); // @[digest.scala 81:19]
  wire [31:0] _GEN_2489 = 6'h37 == state ? $signed(_GEN_1346) : $signed(_GEN_2159); // @[digest.scala 81:19]
  wire [31:0] _GEN_2490 = 6'h37 == state ? $signed(_GEN_1347) : $signed(_GEN_2160); // @[digest.scala 81:19]
  wire [31:0] _GEN_2491 = 6'h37 == state ? $signed(_GEN_1348) : $signed(_GEN_2161); // @[digest.scala 81:19]
  wire [31:0] _GEN_2492 = 6'h37 == state ? $signed(_GEN_1349) : $signed(_GEN_2162); // @[digest.scala 81:19]
  wire [31:0] _GEN_2493 = 6'h37 == state ? $signed(_GEN_1350) : $signed(_GEN_2163); // @[digest.scala 81:19]
  wire [31:0] _GEN_2494 = 6'h37 == state ? $signed(_GEN_1351) : $signed(_GEN_2164); // @[digest.scala 81:19]
  wire [31:0] _GEN_2495 = 6'h37 == state ? $signed(_GEN_1352) : $signed(_GEN_2165); // @[digest.scala 81:19]
  wire [31:0] _GEN_2496 = 6'h37 == state ? $signed(_GEN_1353) : $signed(_GEN_2166); // @[digest.scala 81:19]
  wire [31:0] _GEN_2497 = 6'h37 == state ? $signed(_GEN_1354) : $signed(_GEN_2167); // @[digest.scala 81:19]
  wire [31:0] _GEN_2498 = 6'h37 == state ? $signed(_GEN_1355) : $signed(_GEN_2168); // @[digest.scala 81:19]
  wire [31:0] _GEN_2499 = 6'h37 == state ? $signed(_GEN_1356) : $signed(_GEN_2169); // @[digest.scala 81:19]
  wire [31:0] _GEN_2500 = 6'h37 == state ? $signed(_GEN_1357) : $signed(_GEN_2170); // @[digest.scala 81:19]
  wire [31:0] _GEN_2501 = 6'h37 == state ? $signed(_GEN_1358) : $signed(_GEN_2171); // @[digest.scala 81:19]
  wire [31:0] _GEN_2502 = 6'h37 == state ? $signed(_GEN_1359) : $signed(_GEN_2172); // @[digest.scala 81:19]
  wire [31:0] _GEN_2503 = 6'h37 == state ? $signed(_GEN_1360) : $signed(_GEN_2173); // @[digest.scala 81:19]
  wire  _GEN_2505 = 6'h37 == state & __m_fill_1_io_valid_T; // @[digest.scala 81:19 320:33 63:25]
  wire [5:0] _GEN_2506 = 6'h37 == state ? _state_T_19 : _GEN_2176; // @[digest.scala 321:19 81:19]
  wire  _GEN_2589 = 6'h37 == state ? 1'h0 : _GEN_2175; // @[digest.scala 81:19 68:25]
  wire  _GEN_2672 = 6'h37 == state ? 1'h0 : _GEN_2259; // @[digest.scala 81:19 73:25]
  wire  _GEN_2755 = 6'h37 == state ? 1'h0 : _GEN_2342; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_2837 = 6'h36 == state ? $signed(_GEN_1201) : $signed(_GEN_2424); // @[digest.scala 81:19]
  wire [31:0] _GEN_2838 = 6'h36 == state ? $signed(_GEN_1202) : $signed(_GEN_2425); // @[digest.scala 81:19]
  wire [31:0] _GEN_2839 = 6'h36 == state ? $signed(_GEN_1203) : $signed(_GEN_2426); // @[digest.scala 81:19]
  wire [31:0] _GEN_2840 = 6'h36 == state ? $signed(_GEN_1204) : $signed(_GEN_2427); // @[digest.scala 81:19]
  wire [31:0] _GEN_2841 = 6'h36 == state ? $signed(_GEN_1205) : $signed(_GEN_2428); // @[digest.scala 81:19]
  wire [31:0] _GEN_2842 = 6'h36 == state ? $signed(_GEN_1206) : $signed(_GEN_2429); // @[digest.scala 81:19]
  wire [31:0] _GEN_2843 = 6'h36 == state ? $signed(_GEN_1207) : $signed(_GEN_2430); // @[digest.scala 81:19]
  wire [31:0] _GEN_2844 = 6'h36 == state ? $signed(_GEN_1208) : $signed(_GEN_2431); // @[digest.scala 81:19]
  wire [31:0] _GEN_2845 = 6'h36 == state ? $signed(_GEN_1209) : $signed(_GEN_2432); // @[digest.scala 81:19]
  wire [31:0] _GEN_2846 = 6'h36 == state ? $signed(_GEN_1210) : $signed(_GEN_2433); // @[digest.scala 81:19]
  wire [31:0] _GEN_2847 = 6'h36 == state ? $signed(_GEN_1211) : $signed(_GEN_2434); // @[digest.scala 81:19]
  wire [31:0] _GEN_2848 = 6'h36 == state ? $signed(_GEN_1212) : $signed(_GEN_2435); // @[digest.scala 81:19]
  wire [31:0] _GEN_2849 = 6'h36 == state ? $signed(_GEN_1213) : $signed(_GEN_2436); // @[digest.scala 81:19]
  wire [31:0] _GEN_2850 = 6'h36 == state ? $signed(_GEN_1214) : $signed(_GEN_2437); // @[digest.scala 81:19]
  wire [31:0] _GEN_2851 = 6'h36 == state ? $signed(_GEN_1215) : $signed(_GEN_2438); // @[digest.scala 81:19]
  wire [31:0] _GEN_2852 = 6'h36 == state ? $signed(_GEN_1216) : $signed(_GEN_2439); // @[digest.scala 81:19]
  wire [31:0] _GEN_2853 = 6'h36 == state ? $signed(_GEN_1217) : $signed(_GEN_2440); // @[digest.scala 81:19]
  wire [31:0] _GEN_2854 = 6'h36 == state ? $signed(_GEN_1218) : $signed(_GEN_2441); // @[digest.scala 81:19]
  wire [31:0] _GEN_2855 = 6'h36 == state ? $signed(_GEN_1219) : $signed(_GEN_2442); // @[digest.scala 81:19]
  wire [31:0] _GEN_2856 = 6'h36 == state ? $signed(_GEN_1220) : $signed(_GEN_2443); // @[digest.scala 81:19]
  wire [31:0] _GEN_2857 = 6'h36 == state ? $signed(_GEN_1221) : $signed(_GEN_2444); // @[digest.scala 81:19]
  wire [31:0] _GEN_2858 = 6'h36 == state ? $signed(_GEN_1222) : $signed(_GEN_2445); // @[digest.scala 81:19]
  wire [31:0] _GEN_2859 = 6'h36 == state ? $signed(_GEN_1223) : $signed(_GEN_2446); // @[digest.scala 81:19]
  wire [31:0] _GEN_2860 = 6'h36 == state ? $signed(_GEN_1224) : $signed(_GEN_2447); // @[digest.scala 81:19]
  wire [31:0] _GEN_2861 = 6'h36 == state ? $signed(_GEN_1225) : $signed(_GEN_2448); // @[digest.scala 81:19]
  wire [31:0] _GEN_2862 = 6'h36 == state ? $signed(_GEN_1226) : $signed(_GEN_2449); // @[digest.scala 81:19]
  wire [31:0] _GEN_2863 = 6'h36 == state ? $signed(_GEN_1227) : $signed(_GEN_2450); // @[digest.scala 81:19]
  wire [31:0] _GEN_2864 = 6'h36 == state ? $signed(_GEN_1228) : $signed(_GEN_2451); // @[digest.scala 81:19]
  wire [31:0] _GEN_2865 = 6'h36 == state ? $signed(_GEN_1229) : $signed(_GEN_2452); // @[digest.scala 81:19]
  wire [31:0] _GEN_2866 = 6'h36 == state ? $signed(_GEN_1230) : $signed(_GEN_2453); // @[digest.scala 81:19]
  wire [31:0] _GEN_2867 = 6'h36 == state ? $signed(_GEN_1231) : $signed(_GEN_2454); // @[digest.scala 81:19]
  wire [31:0] _GEN_2868 = 6'h36 == state ? $signed(_GEN_1232) : $signed(_GEN_2455); // @[digest.scala 81:19]
  wire [31:0] _GEN_2869 = 6'h36 == state ? $signed(_GEN_1233) : $signed(_GEN_2456); // @[digest.scala 81:19]
  wire [31:0] _GEN_2870 = 6'h36 == state ? $signed(_GEN_1234) : $signed(_GEN_2457); // @[digest.scala 81:19]
  wire [31:0] _GEN_2871 = 6'h36 == state ? $signed(_GEN_1235) : $signed(_GEN_2458); // @[digest.scala 81:19]
  wire [31:0] _GEN_2872 = 6'h36 == state ? $signed(_GEN_1236) : $signed(_GEN_2459); // @[digest.scala 81:19]
  wire [31:0] _GEN_2873 = 6'h36 == state ? $signed(_GEN_1237) : $signed(_GEN_2460); // @[digest.scala 81:19]
  wire [31:0] _GEN_2874 = 6'h36 == state ? $signed(_GEN_1238) : $signed(_GEN_2461); // @[digest.scala 81:19]
  wire [31:0] _GEN_2875 = 6'h36 == state ? $signed(_GEN_1239) : $signed(_GEN_2462); // @[digest.scala 81:19]
  wire [31:0] _GEN_2876 = 6'h36 == state ? $signed(_GEN_1240) : $signed(_GEN_2463); // @[digest.scala 81:19]
  wire [31:0] _GEN_2877 = 6'h36 == state ? $signed(_GEN_1241) : $signed(_GEN_2464); // @[digest.scala 81:19]
  wire [31:0] _GEN_2878 = 6'h36 == state ? $signed(_GEN_1242) : $signed(_GEN_2465); // @[digest.scala 81:19]
  wire [31:0] _GEN_2879 = 6'h36 == state ? $signed(_GEN_1243) : $signed(_GEN_2466); // @[digest.scala 81:19]
  wire [31:0] _GEN_2880 = 6'h36 == state ? $signed(_GEN_1244) : $signed(_GEN_2467); // @[digest.scala 81:19]
  wire [31:0] _GEN_2881 = 6'h36 == state ? $signed(_GEN_1245) : $signed(_GEN_2468); // @[digest.scala 81:19]
  wire [31:0] _GEN_2882 = 6'h36 == state ? $signed(_GEN_1246) : $signed(_GEN_2469); // @[digest.scala 81:19]
  wire [31:0] _GEN_2883 = 6'h36 == state ? $signed(_GEN_1247) : $signed(_GEN_2470); // @[digest.scala 81:19]
  wire [31:0] _GEN_2884 = 6'h36 == state ? $signed(_GEN_1248) : $signed(_GEN_2471); // @[digest.scala 81:19]
  wire [31:0] _GEN_2885 = 6'h36 == state ? $signed(_GEN_1249) : $signed(_GEN_2472); // @[digest.scala 81:19]
  wire [31:0] _GEN_2886 = 6'h36 == state ? $signed(_GEN_1250) : $signed(_GEN_2473); // @[digest.scala 81:19]
  wire [31:0] _GEN_2887 = 6'h36 == state ? $signed(_GEN_1251) : $signed(_GEN_2474); // @[digest.scala 81:19]
  wire [31:0] _GEN_2888 = 6'h36 == state ? $signed(_GEN_1252) : $signed(_GEN_2475); // @[digest.scala 81:19]
  wire [31:0] _GEN_2889 = 6'h36 == state ? $signed(_GEN_1253) : $signed(_GEN_2476); // @[digest.scala 81:19]
  wire [31:0] _GEN_2890 = 6'h36 == state ? $signed(_GEN_1254) : $signed(_GEN_2477); // @[digest.scala 81:19]
  wire [31:0] _GEN_2891 = 6'h36 == state ? $signed(_GEN_1255) : $signed(_GEN_2478); // @[digest.scala 81:19]
  wire [31:0] _GEN_2892 = 6'h36 == state ? $signed(_GEN_1256) : $signed(_GEN_2479); // @[digest.scala 81:19]
  wire [31:0] _GEN_2893 = 6'h36 == state ? $signed(_GEN_1257) : $signed(_GEN_2480); // @[digest.scala 81:19]
  wire [31:0] _GEN_2894 = 6'h36 == state ? $signed(_GEN_1258) : $signed(_GEN_2481); // @[digest.scala 81:19]
  wire [31:0] _GEN_2895 = 6'h36 == state ? $signed(_GEN_1259) : $signed(_GEN_2482); // @[digest.scala 81:19]
  wire [31:0] _GEN_2896 = 6'h36 == state ? $signed(_GEN_1260) : $signed(_GEN_2483); // @[digest.scala 81:19]
  wire [31:0] _GEN_2897 = 6'h36 == state ? $signed(_GEN_1261) : $signed(_GEN_2484); // @[digest.scala 81:19]
  wire [31:0] _GEN_2898 = 6'h36 == state ? $signed(_GEN_1262) : $signed(_GEN_2485); // @[digest.scala 81:19]
  wire [31:0] _GEN_2899 = 6'h36 == state ? $signed(_GEN_1263) : $signed(_GEN_2486); // @[digest.scala 81:19]
  wire [31:0] _GEN_2900 = 6'h36 == state ? $signed(_GEN_1264) : $signed(_GEN_2487); // @[digest.scala 81:19]
  wire [31:0] _GEN_2901 = 6'h36 == state ? $signed(_GEN_1265) : $signed(_GEN_2488); // @[digest.scala 81:19]
  wire [31:0] _GEN_2902 = 6'h36 == state ? $signed(_GEN_1266) : $signed(_GEN_2489); // @[digest.scala 81:19]
  wire [31:0] _GEN_2903 = 6'h36 == state ? $signed(_GEN_1267) : $signed(_GEN_2490); // @[digest.scala 81:19]
  wire [31:0] _GEN_2904 = 6'h36 == state ? $signed(_GEN_1268) : $signed(_GEN_2491); // @[digest.scala 81:19]
  wire [31:0] _GEN_2905 = 6'h36 == state ? $signed(_GEN_1269) : $signed(_GEN_2492); // @[digest.scala 81:19]
  wire [31:0] _GEN_2906 = 6'h36 == state ? $signed(_GEN_1270) : $signed(_GEN_2493); // @[digest.scala 81:19]
  wire [31:0] _GEN_2907 = 6'h36 == state ? $signed(_GEN_1271) : $signed(_GEN_2494); // @[digest.scala 81:19]
  wire [31:0] _GEN_2908 = 6'h36 == state ? $signed(_GEN_1272) : $signed(_GEN_2495); // @[digest.scala 81:19]
  wire [31:0] _GEN_2909 = 6'h36 == state ? $signed(_GEN_1273) : $signed(_GEN_2496); // @[digest.scala 81:19]
  wire [31:0] _GEN_2910 = 6'h36 == state ? $signed(_GEN_1274) : $signed(_GEN_2497); // @[digest.scala 81:19]
  wire [31:0] _GEN_2911 = 6'h36 == state ? $signed(_GEN_1275) : $signed(_GEN_2498); // @[digest.scala 81:19]
  wire [31:0] _GEN_2912 = 6'h36 == state ? $signed(_GEN_1276) : $signed(_GEN_2499); // @[digest.scala 81:19]
  wire [31:0] _GEN_2913 = 6'h36 == state ? $signed(_GEN_1277) : $signed(_GEN_2500); // @[digest.scala 81:19]
  wire [31:0] _GEN_2914 = 6'h36 == state ? $signed(_GEN_1278) : $signed(_GEN_2501); // @[digest.scala 81:19]
  wire [31:0] _GEN_2915 = 6'h36 == state ? $signed(_GEN_1279) : $signed(_GEN_2502); // @[digest.scala 81:19]
  wire [31:0] _GEN_2916 = 6'h36 == state ? $signed(_GEN_1280) : $signed(_GEN_2503); // @[digest.scala 81:19]
  wire  _GEN_2918 = 6'h36 == state & __m_fill_0_io_valid_T; // @[digest.scala 81:19 310:33 58:25]
  wire [5:0] _GEN_2919 = 6'h36 == state ? _state_T_18 : _GEN_2506; // @[digest.scala 311:19 81:19]
  wire  _GEN_3002 = 6'h36 == state ? 1'h0 : _GEN_2505; // @[digest.scala 81:19 63:25]
  wire  _GEN_3085 = 6'h36 == state ? 1'h0 : _GEN_2589; // @[digest.scala 81:19 68:25]
  wire  _GEN_3168 = 6'h36 == state ? 1'h0 : _GEN_2672; // @[digest.scala 81:19 73:25]
  wire  _GEN_3251 = 6'h36 == state ? 1'h0 : _GEN_2755; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_3252 = 6'h35 == state ? $signed(_i_T_5) : $signed(i); // @[digest.scala 300:15 23:16 81:19]
  wire [5:0] _GEN_3253 = 6'h35 == state ? 6'h36 : _GEN_2919; // @[digest.scala 301:19 81:19]
  wire [31:0] _GEN_3335 = 6'h35 == state ? $signed(digest_0) : $signed(_GEN_2837); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3336 = 6'h35 == state ? $signed(digest_1) : $signed(_GEN_2838); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3337 = 6'h35 == state ? $signed(digest_2) : $signed(_GEN_2839); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3338 = 6'h35 == state ? $signed(digest_3) : $signed(_GEN_2840); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3339 = 6'h35 == state ? $signed(digest_4) : $signed(_GEN_2841); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3340 = 6'h35 == state ? $signed(digest_5) : $signed(_GEN_2842); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3341 = 6'h35 == state ? $signed(digest_6) : $signed(_GEN_2843); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3342 = 6'h35 == state ? $signed(digest_7) : $signed(_GEN_2844); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3343 = 6'h35 == state ? $signed(digest_8) : $signed(_GEN_2845); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3344 = 6'h35 == state ? $signed(digest_9) : $signed(_GEN_2846); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3345 = 6'h35 == state ? $signed(digest_10) : $signed(_GEN_2847); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3346 = 6'h35 == state ? $signed(digest_11) : $signed(_GEN_2848); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3347 = 6'h35 == state ? $signed(digest_12) : $signed(_GEN_2849); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3348 = 6'h35 == state ? $signed(digest_13) : $signed(_GEN_2850); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3349 = 6'h35 == state ? $signed(digest_14) : $signed(_GEN_2851); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3350 = 6'h35 == state ? $signed(digest_15) : $signed(_GEN_2852); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3351 = 6'h35 == state ? $signed(digest_16) : $signed(_GEN_2853); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3352 = 6'h35 == state ? $signed(digest_17) : $signed(_GEN_2854); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3353 = 6'h35 == state ? $signed(digest_18) : $signed(_GEN_2855); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3354 = 6'h35 == state ? $signed(digest_19) : $signed(_GEN_2856); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3355 = 6'h35 == state ? $signed(digest_20) : $signed(_GEN_2857); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3356 = 6'h35 == state ? $signed(digest_21) : $signed(_GEN_2858); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3357 = 6'h35 == state ? $signed(digest_22) : $signed(_GEN_2859); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3358 = 6'h35 == state ? $signed(digest_23) : $signed(_GEN_2860); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3359 = 6'h35 == state ? $signed(digest_24) : $signed(_GEN_2861); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3360 = 6'h35 == state ? $signed(digest_25) : $signed(_GEN_2862); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3361 = 6'h35 == state ? $signed(digest_26) : $signed(_GEN_2863); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3362 = 6'h35 == state ? $signed(digest_27) : $signed(_GEN_2864); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3363 = 6'h35 == state ? $signed(digest_28) : $signed(_GEN_2865); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3364 = 6'h35 == state ? $signed(digest_29) : $signed(_GEN_2866); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3365 = 6'h35 == state ? $signed(digest_30) : $signed(_GEN_2867); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3366 = 6'h35 == state ? $signed(digest_31) : $signed(_GEN_2868); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3367 = 6'h35 == state ? $signed(digest_32) : $signed(_GEN_2869); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3368 = 6'h35 == state ? $signed(digest_33) : $signed(_GEN_2870); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3369 = 6'h35 == state ? $signed(digest_34) : $signed(_GEN_2871); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3370 = 6'h35 == state ? $signed(digest_35) : $signed(_GEN_2872); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3371 = 6'h35 == state ? $signed(digest_36) : $signed(_GEN_2873); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3372 = 6'h35 == state ? $signed(digest_37) : $signed(_GEN_2874); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3373 = 6'h35 == state ? $signed(digest_38) : $signed(_GEN_2875); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3374 = 6'h35 == state ? $signed(digest_39) : $signed(_GEN_2876); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3375 = 6'h35 == state ? $signed(digest_40) : $signed(_GEN_2877); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3376 = 6'h35 == state ? $signed(digest_41) : $signed(_GEN_2878); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3377 = 6'h35 == state ? $signed(digest_42) : $signed(_GEN_2879); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3378 = 6'h35 == state ? $signed(digest_43) : $signed(_GEN_2880); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3379 = 6'h35 == state ? $signed(digest_44) : $signed(_GEN_2881); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3380 = 6'h35 == state ? $signed(digest_45) : $signed(_GEN_2882); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3381 = 6'h35 == state ? $signed(digest_46) : $signed(_GEN_2883); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3382 = 6'h35 == state ? $signed(digest_47) : $signed(_GEN_2884); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3383 = 6'h35 == state ? $signed(digest_48) : $signed(_GEN_2885); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3384 = 6'h35 == state ? $signed(digest_49) : $signed(_GEN_2886); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3385 = 6'h35 == state ? $signed(digest_50) : $signed(_GEN_2887); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3386 = 6'h35 == state ? $signed(digest_51) : $signed(_GEN_2888); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3387 = 6'h35 == state ? $signed(digest_52) : $signed(_GEN_2889); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3388 = 6'h35 == state ? $signed(digest_53) : $signed(_GEN_2890); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3389 = 6'h35 == state ? $signed(digest_54) : $signed(_GEN_2891); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3390 = 6'h35 == state ? $signed(digest_55) : $signed(_GEN_2892); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3391 = 6'h35 == state ? $signed(digest_56) : $signed(_GEN_2893); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3392 = 6'h35 == state ? $signed(digest_57) : $signed(_GEN_2894); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3393 = 6'h35 == state ? $signed(digest_58) : $signed(_GEN_2895); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3394 = 6'h35 == state ? $signed(digest_59) : $signed(_GEN_2896); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3395 = 6'h35 == state ? $signed(digest_60) : $signed(_GEN_2897); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3396 = 6'h35 == state ? $signed(digest_61) : $signed(_GEN_2898); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3397 = 6'h35 == state ? $signed(digest_62) : $signed(_GEN_2899); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3398 = 6'h35 == state ? $signed(digest_63) : $signed(_GEN_2900); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3399 = 6'h35 == state ? $signed(digest_64) : $signed(_GEN_2901); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3400 = 6'h35 == state ? $signed(digest_65) : $signed(_GEN_2902); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3401 = 6'h35 == state ? $signed(digest_66) : $signed(_GEN_2903); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3402 = 6'h35 == state ? $signed(digest_67) : $signed(_GEN_2904); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3403 = 6'h35 == state ? $signed(digest_68) : $signed(_GEN_2905); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3404 = 6'h35 == state ? $signed(digest_69) : $signed(_GEN_2906); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3405 = 6'h35 == state ? $signed(digest_70) : $signed(_GEN_2907); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3406 = 6'h35 == state ? $signed(digest_71) : $signed(_GEN_2908); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3407 = 6'h35 == state ? $signed(digest_72) : $signed(_GEN_2909); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3408 = 6'h35 == state ? $signed(digest_73) : $signed(_GEN_2910); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3409 = 6'h35 == state ? $signed(digest_74) : $signed(_GEN_2911); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3410 = 6'h35 == state ? $signed(digest_75) : $signed(_GEN_2912); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3411 = 6'h35 == state ? $signed(digest_76) : $signed(_GEN_2913); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3412 = 6'h35 == state ? $signed(digest_77) : $signed(_GEN_2914); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3413 = 6'h35 == state ? $signed(digest_78) : $signed(_GEN_2915); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3414 = 6'h35 == state ? $signed(digest_79) : $signed(_GEN_2916); // @[digest.scala 81:19 53:21]
  wire  _GEN_3416 = 6'h35 == state ? 1'h0 : _GEN_2918; // @[digest.scala 81:19 58:25]
  wire  _GEN_3499 = 6'h35 == state ? 1'h0 : _GEN_3002; // @[digest.scala 81:19 63:25]
  wire  _GEN_3582 = 6'h35 == state ? 1'h0 : _GEN_3085; // @[digest.scala 81:19 68:25]
  wire  _GEN_3665 = 6'h35 == state ? 1'h0 : _GEN_3168; // @[digest.scala 81:19 73:25]
  wire  _GEN_3748 = 6'h35 == state ? 1'h0 : _GEN_3251; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_3749 = 6'h34 == state ? $signed(_e_T_2) : $signed(e); // @[digest.scala 296:15 28:16 81:19]
  wire [5:0] _GEN_3750 = 6'h34 == state ? 6'h35 : _GEN_3253; // @[digest.scala 297:19 81:19]
  wire [31:0] _GEN_3751 = 6'h34 == state ? $signed(i) : $signed(_GEN_3252); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_3833 = 6'h34 == state ? $signed(digest_0) : $signed(_GEN_3335); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3834 = 6'h34 == state ? $signed(digest_1) : $signed(_GEN_3336); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3835 = 6'h34 == state ? $signed(digest_2) : $signed(_GEN_3337); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3836 = 6'h34 == state ? $signed(digest_3) : $signed(_GEN_3338); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3837 = 6'h34 == state ? $signed(digest_4) : $signed(_GEN_3339); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3838 = 6'h34 == state ? $signed(digest_5) : $signed(_GEN_3340); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3839 = 6'h34 == state ? $signed(digest_6) : $signed(_GEN_3341); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3840 = 6'h34 == state ? $signed(digest_7) : $signed(_GEN_3342); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3841 = 6'h34 == state ? $signed(digest_8) : $signed(_GEN_3343); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3842 = 6'h34 == state ? $signed(digest_9) : $signed(_GEN_3344); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3843 = 6'h34 == state ? $signed(digest_10) : $signed(_GEN_3345); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3844 = 6'h34 == state ? $signed(digest_11) : $signed(_GEN_3346); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3845 = 6'h34 == state ? $signed(digest_12) : $signed(_GEN_3347); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3846 = 6'h34 == state ? $signed(digest_13) : $signed(_GEN_3348); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3847 = 6'h34 == state ? $signed(digest_14) : $signed(_GEN_3349); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3848 = 6'h34 == state ? $signed(digest_15) : $signed(_GEN_3350); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3849 = 6'h34 == state ? $signed(digest_16) : $signed(_GEN_3351); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3850 = 6'h34 == state ? $signed(digest_17) : $signed(_GEN_3352); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3851 = 6'h34 == state ? $signed(digest_18) : $signed(_GEN_3353); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3852 = 6'h34 == state ? $signed(digest_19) : $signed(_GEN_3354); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3853 = 6'h34 == state ? $signed(digest_20) : $signed(_GEN_3355); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3854 = 6'h34 == state ? $signed(digest_21) : $signed(_GEN_3356); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3855 = 6'h34 == state ? $signed(digest_22) : $signed(_GEN_3357); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3856 = 6'h34 == state ? $signed(digest_23) : $signed(_GEN_3358); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3857 = 6'h34 == state ? $signed(digest_24) : $signed(_GEN_3359); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3858 = 6'h34 == state ? $signed(digest_25) : $signed(_GEN_3360); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3859 = 6'h34 == state ? $signed(digest_26) : $signed(_GEN_3361); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3860 = 6'h34 == state ? $signed(digest_27) : $signed(_GEN_3362); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3861 = 6'h34 == state ? $signed(digest_28) : $signed(_GEN_3363); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3862 = 6'h34 == state ? $signed(digest_29) : $signed(_GEN_3364); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3863 = 6'h34 == state ? $signed(digest_30) : $signed(_GEN_3365); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3864 = 6'h34 == state ? $signed(digest_31) : $signed(_GEN_3366); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3865 = 6'h34 == state ? $signed(digest_32) : $signed(_GEN_3367); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3866 = 6'h34 == state ? $signed(digest_33) : $signed(_GEN_3368); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3867 = 6'h34 == state ? $signed(digest_34) : $signed(_GEN_3369); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3868 = 6'h34 == state ? $signed(digest_35) : $signed(_GEN_3370); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3869 = 6'h34 == state ? $signed(digest_36) : $signed(_GEN_3371); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3870 = 6'h34 == state ? $signed(digest_37) : $signed(_GEN_3372); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3871 = 6'h34 == state ? $signed(digest_38) : $signed(_GEN_3373); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3872 = 6'h34 == state ? $signed(digest_39) : $signed(_GEN_3374); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3873 = 6'h34 == state ? $signed(digest_40) : $signed(_GEN_3375); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3874 = 6'h34 == state ? $signed(digest_41) : $signed(_GEN_3376); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3875 = 6'h34 == state ? $signed(digest_42) : $signed(_GEN_3377); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3876 = 6'h34 == state ? $signed(digest_43) : $signed(_GEN_3378); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3877 = 6'h34 == state ? $signed(digest_44) : $signed(_GEN_3379); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3878 = 6'h34 == state ? $signed(digest_45) : $signed(_GEN_3380); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3879 = 6'h34 == state ? $signed(digest_46) : $signed(_GEN_3381); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3880 = 6'h34 == state ? $signed(digest_47) : $signed(_GEN_3382); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3881 = 6'h34 == state ? $signed(digest_48) : $signed(_GEN_3383); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3882 = 6'h34 == state ? $signed(digest_49) : $signed(_GEN_3384); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3883 = 6'h34 == state ? $signed(digest_50) : $signed(_GEN_3385); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3884 = 6'h34 == state ? $signed(digest_51) : $signed(_GEN_3386); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3885 = 6'h34 == state ? $signed(digest_52) : $signed(_GEN_3387); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3886 = 6'h34 == state ? $signed(digest_53) : $signed(_GEN_3388); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3887 = 6'h34 == state ? $signed(digest_54) : $signed(_GEN_3389); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3888 = 6'h34 == state ? $signed(digest_55) : $signed(_GEN_3390); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3889 = 6'h34 == state ? $signed(digest_56) : $signed(_GEN_3391); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3890 = 6'h34 == state ? $signed(digest_57) : $signed(_GEN_3392); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3891 = 6'h34 == state ? $signed(digest_58) : $signed(_GEN_3393); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3892 = 6'h34 == state ? $signed(digest_59) : $signed(_GEN_3394); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3893 = 6'h34 == state ? $signed(digest_60) : $signed(_GEN_3395); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3894 = 6'h34 == state ? $signed(digest_61) : $signed(_GEN_3396); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3895 = 6'h34 == state ? $signed(digest_62) : $signed(_GEN_3397); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3896 = 6'h34 == state ? $signed(digest_63) : $signed(_GEN_3398); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3897 = 6'h34 == state ? $signed(digest_64) : $signed(_GEN_3399); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3898 = 6'h34 == state ? $signed(digest_65) : $signed(_GEN_3400); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3899 = 6'h34 == state ? $signed(digest_66) : $signed(_GEN_3401); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3900 = 6'h34 == state ? $signed(digest_67) : $signed(_GEN_3402); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3901 = 6'h34 == state ? $signed(digest_68) : $signed(_GEN_3403); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3902 = 6'h34 == state ? $signed(digest_69) : $signed(_GEN_3404); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3903 = 6'h34 == state ? $signed(digest_70) : $signed(_GEN_3405); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3904 = 6'h34 == state ? $signed(digest_71) : $signed(_GEN_3406); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3905 = 6'h34 == state ? $signed(digest_72) : $signed(_GEN_3407); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3906 = 6'h34 == state ? $signed(digest_73) : $signed(_GEN_3408); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3907 = 6'h34 == state ? $signed(digest_74) : $signed(_GEN_3409); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3908 = 6'h34 == state ? $signed(digest_75) : $signed(_GEN_3410); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3909 = 6'h34 == state ? $signed(digest_76) : $signed(_GEN_3411); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3910 = 6'h34 == state ? $signed(digest_77) : $signed(_GEN_3412); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3911 = 6'h34 == state ? $signed(digest_78) : $signed(_GEN_3413); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_3912 = 6'h34 == state ? $signed(digest_79) : $signed(_GEN_3414); // @[digest.scala 81:19 53:21]
  wire  _GEN_3914 = 6'h34 == state ? 1'h0 : _GEN_3416; // @[digest.scala 81:19 58:25]
  wire  _GEN_3997 = 6'h34 == state ? 1'h0 : _GEN_3499; // @[digest.scala 81:19 63:25]
  wire  _GEN_4080 = 6'h34 == state ? 1'h0 : _GEN_3582; // @[digest.scala 81:19 68:25]
  wire  _GEN_4163 = 6'h34 == state ? 1'h0 : _GEN_3665; // @[digest.scala 81:19 73:25]
  wire  _GEN_4246 = 6'h34 == state ? 1'h0 : _GEN_3748; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_4247 = 6'h33 == state ? $signed(_d_T_2) : $signed(d); // @[digest.scala 292:15 27:16 81:19]
  wire [5:0] _GEN_4248 = 6'h33 == state ? 6'h34 : _GEN_3750; // @[digest.scala 293:19 81:19]
  wire [31:0] _GEN_4249 = 6'h33 == state ? $signed(e) : $signed(_GEN_3749); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_4250 = 6'h33 == state ? $signed(i) : $signed(_GEN_3751); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_4332 = 6'h33 == state ? $signed(digest_0) : $signed(_GEN_3833); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4333 = 6'h33 == state ? $signed(digest_1) : $signed(_GEN_3834); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4334 = 6'h33 == state ? $signed(digest_2) : $signed(_GEN_3835); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4335 = 6'h33 == state ? $signed(digest_3) : $signed(_GEN_3836); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4336 = 6'h33 == state ? $signed(digest_4) : $signed(_GEN_3837); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4337 = 6'h33 == state ? $signed(digest_5) : $signed(_GEN_3838); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4338 = 6'h33 == state ? $signed(digest_6) : $signed(_GEN_3839); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4339 = 6'h33 == state ? $signed(digest_7) : $signed(_GEN_3840); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4340 = 6'h33 == state ? $signed(digest_8) : $signed(_GEN_3841); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4341 = 6'h33 == state ? $signed(digest_9) : $signed(_GEN_3842); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4342 = 6'h33 == state ? $signed(digest_10) : $signed(_GEN_3843); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4343 = 6'h33 == state ? $signed(digest_11) : $signed(_GEN_3844); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4344 = 6'h33 == state ? $signed(digest_12) : $signed(_GEN_3845); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4345 = 6'h33 == state ? $signed(digest_13) : $signed(_GEN_3846); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4346 = 6'h33 == state ? $signed(digest_14) : $signed(_GEN_3847); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4347 = 6'h33 == state ? $signed(digest_15) : $signed(_GEN_3848); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4348 = 6'h33 == state ? $signed(digest_16) : $signed(_GEN_3849); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4349 = 6'h33 == state ? $signed(digest_17) : $signed(_GEN_3850); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4350 = 6'h33 == state ? $signed(digest_18) : $signed(_GEN_3851); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4351 = 6'h33 == state ? $signed(digest_19) : $signed(_GEN_3852); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4352 = 6'h33 == state ? $signed(digest_20) : $signed(_GEN_3853); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4353 = 6'h33 == state ? $signed(digest_21) : $signed(_GEN_3854); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4354 = 6'h33 == state ? $signed(digest_22) : $signed(_GEN_3855); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4355 = 6'h33 == state ? $signed(digest_23) : $signed(_GEN_3856); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4356 = 6'h33 == state ? $signed(digest_24) : $signed(_GEN_3857); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4357 = 6'h33 == state ? $signed(digest_25) : $signed(_GEN_3858); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4358 = 6'h33 == state ? $signed(digest_26) : $signed(_GEN_3859); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4359 = 6'h33 == state ? $signed(digest_27) : $signed(_GEN_3860); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4360 = 6'h33 == state ? $signed(digest_28) : $signed(_GEN_3861); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4361 = 6'h33 == state ? $signed(digest_29) : $signed(_GEN_3862); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4362 = 6'h33 == state ? $signed(digest_30) : $signed(_GEN_3863); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4363 = 6'h33 == state ? $signed(digest_31) : $signed(_GEN_3864); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4364 = 6'h33 == state ? $signed(digest_32) : $signed(_GEN_3865); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4365 = 6'h33 == state ? $signed(digest_33) : $signed(_GEN_3866); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4366 = 6'h33 == state ? $signed(digest_34) : $signed(_GEN_3867); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4367 = 6'h33 == state ? $signed(digest_35) : $signed(_GEN_3868); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4368 = 6'h33 == state ? $signed(digest_36) : $signed(_GEN_3869); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4369 = 6'h33 == state ? $signed(digest_37) : $signed(_GEN_3870); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4370 = 6'h33 == state ? $signed(digest_38) : $signed(_GEN_3871); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4371 = 6'h33 == state ? $signed(digest_39) : $signed(_GEN_3872); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4372 = 6'h33 == state ? $signed(digest_40) : $signed(_GEN_3873); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4373 = 6'h33 == state ? $signed(digest_41) : $signed(_GEN_3874); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4374 = 6'h33 == state ? $signed(digest_42) : $signed(_GEN_3875); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4375 = 6'h33 == state ? $signed(digest_43) : $signed(_GEN_3876); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4376 = 6'h33 == state ? $signed(digest_44) : $signed(_GEN_3877); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4377 = 6'h33 == state ? $signed(digest_45) : $signed(_GEN_3878); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4378 = 6'h33 == state ? $signed(digest_46) : $signed(_GEN_3879); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4379 = 6'h33 == state ? $signed(digest_47) : $signed(_GEN_3880); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4380 = 6'h33 == state ? $signed(digest_48) : $signed(_GEN_3881); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4381 = 6'h33 == state ? $signed(digest_49) : $signed(_GEN_3882); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4382 = 6'h33 == state ? $signed(digest_50) : $signed(_GEN_3883); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4383 = 6'h33 == state ? $signed(digest_51) : $signed(_GEN_3884); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4384 = 6'h33 == state ? $signed(digest_52) : $signed(_GEN_3885); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4385 = 6'h33 == state ? $signed(digest_53) : $signed(_GEN_3886); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4386 = 6'h33 == state ? $signed(digest_54) : $signed(_GEN_3887); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4387 = 6'h33 == state ? $signed(digest_55) : $signed(_GEN_3888); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4388 = 6'h33 == state ? $signed(digest_56) : $signed(_GEN_3889); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4389 = 6'h33 == state ? $signed(digest_57) : $signed(_GEN_3890); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4390 = 6'h33 == state ? $signed(digest_58) : $signed(_GEN_3891); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4391 = 6'h33 == state ? $signed(digest_59) : $signed(_GEN_3892); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4392 = 6'h33 == state ? $signed(digest_60) : $signed(_GEN_3893); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4393 = 6'h33 == state ? $signed(digest_61) : $signed(_GEN_3894); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4394 = 6'h33 == state ? $signed(digest_62) : $signed(_GEN_3895); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4395 = 6'h33 == state ? $signed(digest_63) : $signed(_GEN_3896); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4396 = 6'h33 == state ? $signed(digest_64) : $signed(_GEN_3897); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4397 = 6'h33 == state ? $signed(digest_65) : $signed(_GEN_3898); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4398 = 6'h33 == state ? $signed(digest_66) : $signed(_GEN_3899); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4399 = 6'h33 == state ? $signed(digest_67) : $signed(_GEN_3900); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4400 = 6'h33 == state ? $signed(digest_68) : $signed(_GEN_3901); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4401 = 6'h33 == state ? $signed(digest_69) : $signed(_GEN_3902); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4402 = 6'h33 == state ? $signed(digest_70) : $signed(_GEN_3903); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4403 = 6'h33 == state ? $signed(digest_71) : $signed(_GEN_3904); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4404 = 6'h33 == state ? $signed(digest_72) : $signed(_GEN_3905); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4405 = 6'h33 == state ? $signed(digest_73) : $signed(_GEN_3906); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4406 = 6'h33 == state ? $signed(digest_74) : $signed(_GEN_3907); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4407 = 6'h33 == state ? $signed(digest_75) : $signed(_GEN_3908); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4408 = 6'h33 == state ? $signed(digest_76) : $signed(_GEN_3909); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4409 = 6'h33 == state ? $signed(digest_77) : $signed(_GEN_3910); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4410 = 6'h33 == state ? $signed(digest_78) : $signed(_GEN_3911); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4411 = 6'h33 == state ? $signed(digest_79) : $signed(_GEN_3912); // @[digest.scala 81:19 53:21]
  wire  _GEN_4413 = 6'h33 == state ? 1'h0 : _GEN_3914; // @[digest.scala 81:19 58:25]
  wire  _GEN_4496 = 6'h33 == state ? 1'h0 : _GEN_3997; // @[digest.scala 81:19 63:25]
  wire  _GEN_4579 = 6'h33 == state ? 1'h0 : _GEN_4080; // @[digest.scala 81:19 68:25]
  wire  _GEN_4662 = 6'h33 == state ? 1'h0 : _GEN_4163; // @[digest.scala 81:19 73:25]
  wire  _GEN_4745 = 6'h33 == state ? 1'h0 : _GEN_4246; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_4746 = 6'h32 == state ? $signed(_c_T_2) : $signed(c); // @[digest.scala 288:15 26:16 81:19]
  wire [5:0] _GEN_4747 = 6'h32 == state ? 6'h33 : _GEN_4248; // @[digest.scala 289:19 81:19]
  wire [31:0] _GEN_4748 = 6'h32 == state ? $signed(d) : $signed(_GEN_4247); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_4749 = 6'h32 == state ? $signed(e) : $signed(_GEN_4249); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_4750 = 6'h32 == state ? $signed(i) : $signed(_GEN_4250); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_4832 = 6'h32 == state ? $signed(digest_0) : $signed(_GEN_4332); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4833 = 6'h32 == state ? $signed(digest_1) : $signed(_GEN_4333); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4834 = 6'h32 == state ? $signed(digest_2) : $signed(_GEN_4334); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4835 = 6'h32 == state ? $signed(digest_3) : $signed(_GEN_4335); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4836 = 6'h32 == state ? $signed(digest_4) : $signed(_GEN_4336); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4837 = 6'h32 == state ? $signed(digest_5) : $signed(_GEN_4337); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4838 = 6'h32 == state ? $signed(digest_6) : $signed(_GEN_4338); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4839 = 6'h32 == state ? $signed(digest_7) : $signed(_GEN_4339); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4840 = 6'h32 == state ? $signed(digest_8) : $signed(_GEN_4340); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4841 = 6'h32 == state ? $signed(digest_9) : $signed(_GEN_4341); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4842 = 6'h32 == state ? $signed(digest_10) : $signed(_GEN_4342); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4843 = 6'h32 == state ? $signed(digest_11) : $signed(_GEN_4343); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4844 = 6'h32 == state ? $signed(digest_12) : $signed(_GEN_4344); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4845 = 6'h32 == state ? $signed(digest_13) : $signed(_GEN_4345); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4846 = 6'h32 == state ? $signed(digest_14) : $signed(_GEN_4346); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4847 = 6'h32 == state ? $signed(digest_15) : $signed(_GEN_4347); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4848 = 6'h32 == state ? $signed(digest_16) : $signed(_GEN_4348); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4849 = 6'h32 == state ? $signed(digest_17) : $signed(_GEN_4349); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4850 = 6'h32 == state ? $signed(digest_18) : $signed(_GEN_4350); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4851 = 6'h32 == state ? $signed(digest_19) : $signed(_GEN_4351); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4852 = 6'h32 == state ? $signed(digest_20) : $signed(_GEN_4352); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4853 = 6'h32 == state ? $signed(digest_21) : $signed(_GEN_4353); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4854 = 6'h32 == state ? $signed(digest_22) : $signed(_GEN_4354); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4855 = 6'h32 == state ? $signed(digest_23) : $signed(_GEN_4355); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4856 = 6'h32 == state ? $signed(digest_24) : $signed(_GEN_4356); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4857 = 6'h32 == state ? $signed(digest_25) : $signed(_GEN_4357); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4858 = 6'h32 == state ? $signed(digest_26) : $signed(_GEN_4358); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4859 = 6'h32 == state ? $signed(digest_27) : $signed(_GEN_4359); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4860 = 6'h32 == state ? $signed(digest_28) : $signed(_GEN_4360); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4861 = 6'h32 == state ? $signed(digest_29) : $signed(_GEN_4361); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4862 = 6'h32 == state ? $signed(digest_30) : $signed(_GEN_4362); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4863 = 6'h32 == state ? $signed(digest_31) : $signed(_GEN_4363); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4864 = 6'h32 == state ? $signed(digest_32) : $signed(_GEN_4364); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4865 = 6'h32 == state ? $signed(digest_33) : $signed(_GEN_4365); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4866 = 6'h32 == state ? $signed(digest_34) : $signed(_GEN_4366); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4867 = 6'h32 == state ? $signed(digest_35) : $signed(_GEN_4367); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4868 = 6'h32 == state ? $signed(digest_36) : $signed(_GEN_4368); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4869 = 6'h32 == state ? $signed(digest_37) : $signed(_GEN_4369); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4870 = 6'h32 == state ? $signed(digest_38) : $signed(_GEN_4370); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4871 = 6'h32 == state ? $signed(digest_39) : $signed(_GEN_4371); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4872 = 6'h32 == state ? $signed(digest_40) : $signed(_GEN_4372); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4873 = 6'h32 == state ? $signed(digest_41) : $signed(_GEN_4373); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4874 = 6'h32 == state ? $signed(digest_42) : $signed(_GEN_4374); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4875 = 6'h32 == state ? $signed(digest_43) : $signed(_GEN_4375); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4876 = 6'h32 == state ? $signed(digest_44) : $signed(_GEN_4376); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4877 = 6'h32 == state ? $signed(digest_45) : $signed(_GEN_4377); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4878 = 6'h32 == state ? $signed(digest_46) : $signed(_GEN_4378); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4879 = 6'h32 == state ? $signed(digest_47) : $signed(_GEN_4379); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4880 = 6'h32 == state ? $signed(digest_48) : $signed(_GEN_4380); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4881 = 6'h32 == state ? $signed(digest_49) : $signed(_GEN_4381); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4882 = 6'h32 == state ? $signed(digest_50) : $signed(_GEN_4382); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4883 = 6'h32 == state ? $signed(digest_51) : $signed(_GEN_4383); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4884 = 6'h32 == state ? $signed(digest_52) : $signed(_GEN_4384); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4885 = 6'h32 == state ? $signed(digest_53) : $signed(_GEN_4385); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4886 = 6'h32 == state ? $signed(digest_54) : $signed(_GEN_4386); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4887 = 6'h32 == state ? $signed(digest_55) : $signed(_GEN_4387); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4888 = 6'h32 == state ? $signed(digest_56) : $signed(_GEN_4388); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4889 = 6'h32 == state ? $signed(digest_57) : $signed(_GEN_4389); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4890 = 6'h32 == state ? $signed(digest_58) : $signed(_GEN_4390); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4891 = 6'h32 == state ? $signed(digest_59) : $signed(_GEN_4391); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4892 = 6'h32 == state ? $signed(digest_60) : $signed(_GEN_4392); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4893 = 6'h32 == state ? $signed(digest_61) : $signed(_GEN_4393); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4894 = 6'h32 == state ? $signed(digest_62) : $signed(_GEN_4394); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4895 = 6'h32 == state ? $signed(digest_63) : $signed(_GEN_4395); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4896 = 6'h32 == state ? $signed(digest_64) : $signed(_GEN_4396); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4897 = 6'h32 == state ? $signed(digest_65) : $signed(_GEN_4397); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4898 = 6'h32 == state ? $signed(digest_66) : $signed(_GEN_4398); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4899 = 6'h32 == state ? $signed(digest_67) : $signed(_GEN_4399); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4900 = 6'h32 == state ? $signed(digest_68) : $signed(_GEN_4400); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4901 = 6'h32 == state ? $signed(digest_69) : $signed(_GEN_4401); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4902 = 6'h32 == state ? $signed(digest_70) : $signed(_GEN_4402); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4903 = 6'h32 == state ? $signed(digest_71) : $signed(_GEN_4403); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4904 = 6'h32 == state ? $signed(digest_72) : $signed(_GEN_4404); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4905 = 6'h32 == state ? $signed(digest_73) : $signed(_GEN_4405); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4906 = 6'h32 == state ? $signed(digest_74) : $signed(_GEN_4406); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4907 = 6'h32 == state ? $signed(digest_75) : $signed(_GEN_4407); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4908 = 6'h32 == state ? $signed(digest_76) : $signed(_GEN_4408); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4909 = 6'h32 == state ? $signed(digest_77) : $signed(_GEN_4409); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4910 = 6'h32 == state ? $signed(digest_78) : $signed(_GEN_4410); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_4911 = 6'h32 == state ? $signed(digest_79) : $signed(_GEN_4411); // @[digest.scala 81:19 53:21]
  wire  _GEN_4913 = 6'h32 == state ? 1'h0 : _GEN_4413; // @[digest.scala 81:19 58:25]
  wire  _GEN_4996 = 6'h32 == state ? 1'h0 : _GEN_4496; // @[digest.scala 81:19 63:25]
  wire  _GEN_5079 = 6'h32 == state ? 1'h0 : _GEN_4579; // @[digest.scala 81:19 68:25]
  wire  _GEN_5162 = 6'h32 == state ? 1'h0 : _GEN_4662; // @[digest.scala 81:19 73:25]
  wire  _GEN_5245 = 6'h32 == state ? 1'h0 : _GEN_4745; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_5246 = 6'h31 == state ? $signed(_b_T_2) : $signed(b); // @[digest.scala 284:15 25:16 81:19]
  wire [5:0] _GEN_5247 = 6'h31 == state ? 6'h32 : _GEN_4747; // @[digest.scala 285:19 81:19]
  wire [31:0] _GEN_5248 = 6'h31 == state ? $signed(c) : $signed(_GEN_4746); // @[digest.scala 26:16 81:19]
  wire [31:0] _GEN_5249 = 6'h31 == state ? $signed(d) : $signed(_GEN_4748); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_5250 = 6'h31 == state ? $signed(e) : $signed(_GEN_4749); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_5251 = 6'h31 == state ? $signed(i) : $signed(_GEN_4750); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_5333 = 6'h31 == state ? $signed(digest_0) : $signed(_GEN_4832); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5334 = 6'h31 == state ? $signed(digest_1) : $signed(_GEN_4833); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5335 = 6'h31 == state ? $signed(digest_2) : $signed(_GEN_4834); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5336 = 6'h31 == state ? $signed(digest_3) : $signed(_GEN_4835); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5337 = 6'h31 == state ? $signed(digest_4) : $signed(_GEN_4836); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5338 = 6'h31 == state ? $signed(digest_5) : $signed(_GEN_4837); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5339 = 6'h31 == state ? $signed(digest_6) : $signed(_GEN_4838); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5340 = 6'h31 == state ? $signed(digest_7) : $signed(_GEN_4839); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5341 = 6'h31 == state ? $signed(digest_8) : $signed(_GEN_4840); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5342 = 6'h31 == state ? $signed(digest_9) : $signed(_GEN_4841); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5343 = 6'h31 == state ? $signed(digest_10) : $signed(_GEN_4842); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5344 = 6'h31 == state ? $signed(digest_11) : $signed(_GEN_4843); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5345 = 6'h31 == state ? $signed(digest_12) : $signed(_GEN_4844); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5346 = 6'h31 == state ? $signed(digest_13) : $signed(_GEN_4845); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5347 = 6'h31 == state ? $signed(digest_14) : $signed(_GEN_4846); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5348 = 6'h31 == state ? $signed(digest_15) : $signed(_GEN_4847); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5349 = 6'h31 == state ? $signed(digest_16) : $signed(_GEN_4848); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5350 = 6'h31 == state ? $signed(digest_17) : $signed(_GEN_4849); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5351 = 6'h31 == state ? $signed(digest_18) : $signed(_GEN_4850); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5352 = 6'h31 == state ? $signed(digest_19) : $signed(_GEN_4851); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5353 = 6'h31 == state ? $signed(digest_20) : $signed(_GEN_4852); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5354 = 6'h31 == state ? $signed(digest_21) : $signed(_GEN_4853); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5355 = 6'h31 == state ? $signed(digest_22) : $signed(_GEN_4854); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5356 = 6'h31 == state ? $signed(digest_23) : $signed(_GEN_4855); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5357 = 6'h31 == state ? $signed(digest_24) : $signed(_GEN_4856); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5358 = 6'h31 == state ? $signed(digest_25) : $signed(_GEN_4857); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5359 = 6'h31 == state ? $signed(digest_26) : $signed(_GEN_4858); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5360 = 6'h31 == state ? $signed(digest_27) : $signed(_GEN_4859); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5361 = 6'h31 == state ? $signed(digest_28) : $signed(_GEN_4860); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5362 = 6'h31 == state ? $signed(digest_29) : $signed(_GEN_4861); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5363 = 6'h31 == state ? $signed(digest_30) : $signed(_GEN_4862); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5364 = 6'h31 == state ? $signed(digest_31) : $signed(_GEN_4863); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5365 = 6'h31 == state ? $signed(digest_32) : $signed(_GEN_4864); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5366 = 6'h31 == state ? $signed(digest_33) : $signed(_GEN_4865); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5367 = 6'h31 == state ? $signed(digest_34) : $signed(_GEN_4866); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5368 = 6'h31 == state ? $signed(digest_35) : $signed(_GEN_4867); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5369 = 6'h31 == state ? $signed(digest_36) : $signed(_GEN_4868); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5370 = 6'h31 == state ? $signed(digest_37) : $signed(_GEN_4869); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5371 = 6'h31 == state ? $signed(digest_38) : $signed(_GEN_4870); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5372 = 6'h31 == state ? $signed(digest_39) : $signed(_GEN_4871); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5373 = 6'h31 == state ? $signed(digest_40) : $signed(_GEN_4872); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5374 = 6'h31 == state ? $signed(digest_41) : $signed(_GEN_4873); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5375 = 6'h31 == state ? $signed(digest_42) : $signed(_GEN_4874); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5376 = 6'h31 == state ? $signed(digest_43) : $signed(_GEN_4875); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5377 = 6'h31 == state ? $signed(digest_44) : $signed(_GEN_4876); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5378 = 6'h31 == state ? $signed(digest_45) : $signed(_GEN_4877); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5379 = 6'h31 == state ? $signed(digest_46) : $signed(_GEN_4878); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5380 = 6'h31 == state ? $signed(digest_47) : $signed(_GEN_4879); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5381 = 6'h31 == state ? $signed(digest_48) : $signed(_GEN_4880); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5382 = 6'h31 == state ? $signed(digest_49) : $signed(_GEN_4881); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5383 = 6'h31 == state ? $signed(digest_50) : $signed(_GEN_4882); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5384 = 6'h31 == state ? $signed(digest_51) : $signed(_GEN_4883); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5385 = 6'h31 == state ? $signed(digest_52) : $signed(_GEN_4884); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5386 = 6'h31 == state ? $signed(digest_53) : $signed(_GEN_4885); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5387 = 6'h31 == state ? $signed(digest_54) : $signed(_GEN_4886); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5388 = 6'h31 == state ? $signed(digest_55) : $signed(_GEN_4887); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5389 = 6'h31 == state ? $signed(digest_56) : $signed(_GEN_4888); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5390 = 6'h31 == state ? $signed(digest_57) : $signed(_GEN_4889); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5391 = 6'h31 == state ? $signed(digest_58) : $signed(_GEN_4890); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5392 = 6'h31 == state ? $signed(digest_59) : $signed(_GEN_4891); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5393 = 6'h31 == state ? $signed(digest_60) : $signed(_GEN_4892); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5394 = 6'h31 == state ? $signed(digest_61) : $signed(_GEN_4893); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5395 = 6'h31 == state ? $signed(digest_62) : $signed(_GEN_4894); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5396 = 6'h31 == state ? $signed(digest_63) : $signed(_GEN_4895); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5397 = 6'h31 == state ? $signed(digest_64) : $signed(_GEN_4896); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5398 = 6'h31 == state ? $signed(digest_65) : $signed(_GEN_4897); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5399 = 6'h31 == state ? $signed(digest_66) : $signed(_GEN_4898); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5400 = 6'h31 == state ? $signed(digest_67) : $signed(_GEN_4899); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5401 = 6'h31 == state ? $signed(digest_68) : $signed(_GEN_4900); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5402 = 6'h31 == state ? $signed(digest_69) : $signed(_GEN_4901); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5403 = 6'h31 == state ? $signed(digest_70) : $signed(_GEN_4902); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5404 = 6'h31 == state ? $signed(digest_71) : $signed(_GEN_4903); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5405 = 6'h31 == state ? $signed(digest_72) : $signed(_GEN_4904); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5406 = 6'h31 == state ? $signed(digest_73) : $signed(_GEN_4905); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5407 = 6'h31 == state ? $signed(digest_74) : $signed(_GEN_4906); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5408 = 6'h31 == state ? $signed(digest_75) : $signed(_GEN_4907); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5409 = 6'h31 == state ? $signed(digest_76) : $signed(_GEN_4908); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5410 = 6'h31 == state ? $signed(digest_77) : $signed(_GEN_4909); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5411 = 6'h31 == state ? $signed(digest_78) : $signed(_GEN_4910); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5412 = 6'h31 == state ? $signed(digest_79) : $signed(_GEN_4911); // @[digest.scala 81:19 53:21]
  wire  _GEN_5414 = 6'h31 == state ? 1'h0 : _GEN_4913; // @[digest.scala 81:19 58:25]
  wire  _GEN_5497 = 6'h31 == state ? 1'h0 : _GEN_4996; // @[digest.scala 81:19 63:25]
  wire  _GEN_5580 = 6'h31 == state ? 1'h0 : _GEN_5079; // @[digest.scala 81:19 68:25]
  wire  _GEN_5663 = 6'h31 == state ? 1'h0 : _GEN_5162; // @[digest.scala 81:19 73:25]
  wire  _GEN_5746 = 6'h31 == state ? 1'h0 : _GEN_5245; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_5747 = 6'h30 == state ? $signed(_a_T_2) : $signed(a); // @[digest.scala 280:15 24:16 81:19]
  wire [5:0] _GEN_5748 = 6'h30 == state ? 6'h31 : _GEN_5247; // @[digest.scala 281:19 81:19]
  wire [31:0] _GEN_5749 = 6'h30 == state ? $signed(b) : $signed(_GEN_5246); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_5750 = 6'h30 == state ? $signed(c) : $signed(_GEN_5248); // @[digest.scala 26:16 81:19]
  wire [31:0] _GEN_5751 = 6'h30 == state ? $signed(d) : $signed(_GEN_5249); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_5752 = 6'h30 == state ? $signed(e) : $signed(_GEN_5250); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_5753 = 6'h30 == state ? $signed(i) : $signed(_GEN_5251); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_5835 = 6'h30 == state ? $signed(digest_0) : $signed(_GEN_5333); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5836 = 6'h30 == state ? $signed(digest_1) : $signed(_GEN_5334); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5837 = 6'h30 == state ? $signed(digest_2) : $signed(_GEN_5335); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5838 = 6'h30 == state ? $signed(digest_3) : $signed(_GEN_5336); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5839 = 6'h30 == state ? $signed(digest_4) : $signed(_GEN_5337); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5840 = 6'h30 == state ? $signed(digest_5) : $signed(_GEN_5338); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5841 = 6'h30 == state ? $signed(digest_6) : $signed(_GEN_5339); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5842 = 6'h30 == state ? $signed(digest_7) : $signed(_GEN_5340); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5843 = 6'h30 == state ? $signed(digest_8) : $signed(_GEN_5341); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5844 = 6'h30 == state ? $signed(digest_9) : $signed(_GEN_5342); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5845 = 6'h30 == state ? $signed(digest_10) : $signed(_GEN_5343); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5846 = 6'h30 == state ? $signed(digest_11) : $signed(_GEN_5344); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5847 = 6'h30 == state ? $signed(digest_12) : $signed(_GEN_5345); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5848 = 6'h30 == state ? $signed(digest_13) : $signed(_GEN_5346); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5849 = 6'h30 == state ? $signed(digest_14) : $signed(_GEN_5347); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5850 = 6'h30 == state ? $signed(digest_15) : $signed(_GEN_5348); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5851 = 6'h30 == state ? $signed(digest_16) : $signed(_GEN_5349); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5852 = 6'h30 == state ? $signed(digest_17) : $signed(_GEN_5350); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5853 = 6'h30 == state ? $signed(digest_18) : $signed(_GEN_5351); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5854 = 6'h30 == state ? $signed(digest_19) : $signed(_GEN_5352); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5855 = 6'h30 == state ? $signed(digest_20) : $signed(_GEN_5353); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5856 = 6'h30 == state ? $signed(digest_21) : $signed(_GEN_5354); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5857 = 6'h30 == state ? $signed(digest_22) : $signed(_GEN_5355); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5858 = 6'h30 == state ? $signed(digest_23) : $signed(_GEN_5356); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5859 = 6'h30 == state ? $signed(digest_24) : $signed(_GEN_5357); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5860 = 6'h30 == state ? $signed(digest_25) : $signed(_GEN_5358); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5861 = 6'h30 == state ? $signed(digest_26) : $signed(_GEN_5359); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5862 = 6'h30 == state ? $signed(digest_27) : $signed(_GEN_5360); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5863 = 6'h30 == state ? $signed(digest_28) : $signed(_GEN_5361); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5864 = 6'h30 == state ? $signed(digest_29) : $signed(_GEN_5362); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5865 = 6'h30 == state ? $signed(digest_30) : $signed(_GEN_5363); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5866 = 6'h30 == state ? $signed(digest_31) : $signed(_GEN_5364); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5867 = 6'h30 == state ? $signed(digest_32) : $signed(_GEN_5365); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5868 = 6'h30 == state ? $signed(digest_33) : $signed(_GEN_5366); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5869 = 6'h30 == state ? $signed(digest_34) : $signed(_GEN_5367); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5870 = 6'h30 == state ? $signed(digest_35) : $signed(_GEN_5368); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5871 = 6'h30 == state ? $signed(digest_36) : $signed(_GEN_5369); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5872 = 6'h30 == state ? $signed(digest_37) : $signed(_GEN_5370); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5873 = 6'h30 == state ? $signed(digest_38) : $signed(_GEN_5371); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5874 = 6'h30 == state ? $signed(digest_39) : $signed(_GEN_5372); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5875 = 6'h30 == state ? $signed(digest_40) : $signed(_GEN_5373); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5876 = 6'h30 == state ? $signed(digest_41) : $signed(_GEN_5374); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5877 = 6'h30 == state ? $signed(digest_42) : $signed(_GEN_5375); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5878 = 6'h30 == state ? $signed(digest_43) : $signed(_GEN_5376); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5879 = 6'h30 == state ? $signed(digest_44) : $signed(_GEN_5377); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5880 = 6'h30 == state ? $signed(digest_45) : $signed(_GEN_5378); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5881 = 6'h30 == state ? $signed(digest_46) : $signed(_GEN_5379); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5882 = 6'h30 == state ? $signed(digest_47) : $signed(_GEN_5380); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5883 = 6'h30 == state ? $signed(digest_48) : $signed(_GEN_5381); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5884 = 6'h30 == state ? $signed(digest_49) : $signed(_GEN_5382); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5885 = 6'h30 == state ? $signed(digest_50) : $signed(_GEN_5383); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5886 = 6'h30 == state ? $signed(digest_51) : $signed(_GEN_5384); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5887 = 6'h30 == state ? $signed(digest_52) : $signed(_GEN_5385); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5888 = 6'h30 == state ? $signed(digest_53) : $signed(_GEN_5386); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5889 = 6'h30 == state ? $signed(digest_54) : $signed(_GEN_5387); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5890 = 6'h30 == state ? $signed(digest_55) : $signed(_GEN_5388); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5891 = 6'h30 == state ? $signed(digest_56) : $signed(_GEN_5389); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5892 = 6'h30 == state ? $signed(digest_57) : $signed(_GEN_5390); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5893 = 6'h30 == state ? $signed(digest_58) : $signed(_GEN_5391); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5894 = 6'h30 == state ? $signed(digest_59) : $signed(_GEN_5392); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5895 = 6'h30 == state ? $signed(digest_60) : $signed(_GEN_5393); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5896 = 6'h30 == state ? $signed(digest_61) : $signed(_GEN_5394); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5897 = 6'h30 == state ? $signed(digest_62) : $signed(_GEN_5395); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5898 = 6'h30 == state ? $signed(digest_63) : $signed(_GEN_5396); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5899 = 6'h30 == state ? $signed(digest_64) : $signed(_GEN_5397); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5900 = 6'h30 == state ? $signed(digest_65) : $signed(_GEN_5398); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5901 = 6'h30 == state ? $signed(digest_66) : $signed(_GEN_5399); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5902 = 6'h30 == state ? $signed(digest_67) : $signed(_GEN_5400); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5903 = 6'h30 == state ? $signed(digest_68) : $signed(_GEN_5401); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5904 = 6'h30 == state ? $signed(digest_69) : $signed(_GEN_5402); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5905 = 6'h30 == state ? $signed(digest_70) : $signed(_GEN_5403); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5906 = 6'h30 == state ? $signed(digest_71) : $signed(_GEN_5404); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5907 = 6'h30 == state ? $signed(digest_72) : $signed(_GEN_5405); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5908 = 6'h30 == state ? $signed(digest_73) : $signed(_GEN_5406); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5909 = 6'h30 == state ? $signed(digest_74) : $signed(_GEN_5407); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5910 = 6'h30 == state ? $signed(digest_75) : $signed(_GEN_5408); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5911 = 6'h30 == state ? $signed(digest_76) : $signed(_GEN_5409); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5912 = 6'h30 == state ? $signed(digest_77) : $signed(_GEN_5410); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5913 = 6'h30 == state ? $signed(digest_78) : $signed(_GEN_5411); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_5914 = 6'h30 == state ? $signed(digest_79) : $signed(_GEN_5412); // @[digest.scala 81:19 53:21]
  wire  _GEN_5916 = 6'h30 == state ? 1'h0 : _GEN_5414; // @[digest.scala 81:19 58:25]
  wire  _GEN_5999 = 6'h30 == state ? 1'h0 : _GEN_5497; // @[digest.scala 81:19 63:25]
  wire  _GEN_6082 = 6'h30 == state ? 1'h0 : _GEN_5580; // @[digest.scala 81:19 68:25]
  wire  _GEN_6165 = 6'h30 == state ? 1'h0 : _GEN_5663; // @[digest.scala 81:19 73:25]
  wire  _GEN_6248 = 6'h30 == state ? 1'h0 : _GEN_5746; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_6249 = 6'h2f == state ? $signed(_j_T_2) : $signed(j); // @[digest.scala 276:15 34:16 81:19]
  wire [5:0] _GEN_6250 = 6'h2f == state ? 6'h17 : _GEN_5748; // @[digest.scala 277:19 81:19]
  wire [31:0] _GEN_6251 = 6'h2f == state ? $signed(a) : $signed(_GEN_5747); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_6252 = 6'h2f == state ? $signed(b) : $signed(_GEN_5749); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_6253 = 6'h2f == state ? $signed(c) : $signed(_GEN_5750); // @[digest.scala 26:16 81:19]
  wire [31:0] _GEN_6254 = 6'h2f == state ? $signed(d) : $signed(_GEN_5751); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_6255 = 6'h2f == state ? $signed(e) : $signed(_GEN_5752); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_6256 = 6'h2f == state ? $signed(i) : $signed(_GEN_5753); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_6338 = 6'h2f == state ? $signed(digest_0) : $signed(_GEN_5835); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6339 = 6'h2f == state ? $signed(digest_1) : $signed(_GEN_5836); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6340 = 6'h2f == state ? $signed(digest_2) : $signed(_GEN_5837); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6341 = 6'h2f == state ? $signed(digest_3) : $signed(_GEN_5838); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6342 = 6'h2f == state ? $signed(digest_4) : $signed(_GEN_5839); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6343 = 6'h2f == state ? $signed(digest_5) : $signed(_GEN_5840); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6344 = 6'h2f == state ? $signed(digest_6) : $signed(_GEN_5841); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6345 = 6'h2f == state ? $signed(digest_7) : $signed(_GEN_5842); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6346 = 6'h2f == state ? $signed(digest_8) : $signed(_GEN_5843); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6347 = 6'h2f == state ? $signed(digest_9) : $signed(_GEN_5844); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6348 = 6'h2f == state ? $signed(digest_10) : $signed(_GEN_5845); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6349 = 6'h2f == state ? $signed(digest_11) : $signed(_GEN_5846); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6350 = 6'h2f == state ? $signed(digest_12) : $signed(_GEN_5847); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6351 = 6'h2f == state ? $signed(digest_13) : $signed(_GEN_5848); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6352 = 6'h2f == state ? $signed(digest_14) : $signed(_GEN_5849); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6353 = 6'h2f == state ? $signed(digest_15) : $signed(_GEN_5850); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6354 = 6'h2f == state ? $signed(digest_16) : $signed(_GEN_5851); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6355 = 6'h2f == state ? $signed(digest_17) : $signed(_GEN_5852); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6356 = 6'h2f == state ? $signed(digest_18) : $signed(_GEN_5853); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6357 = 6'h2f == state ? $signed(digest_19) : $signed(_GEN_5854); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6358 = 6'h2f == state ? $signed(digest_20) : $signed(_GEN_5855); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6359 = 6'h2f == state ? $signed(digest_21) : $signed(_GEN_5856); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6360 = 6'h2f == state ? $signed(digest_22) : $signed(_GEN_5857); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6361 = 6'h2f == state ? $signed(digest_23) : $signed(_GEN_5858); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6362 = 6'h2f == state ? $signed(digest_24) : $signed(_GEN_5859); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6363 = 6'h2f == state ? $signed(digest_25) : $signed(_GEN_5860); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6364 = 6'h2f == state ? $signed(digest_26) : $signed(_GEN_5861); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6365 = 6'h2f == state ? $signed(digest_27) : $signed(_GEN_5862); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6366 = 6'h2f == state ? $signed(digest_28) : $signed(_GEN_5863); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6367 = 6'h2f == state ? $signed(digest_29) : $signed(_GEN_5864); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6368 = 6'h2f == state ? $signed(digest_30) : $signed(_GEN_5865); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6369 = 6'h2f == state ? $signed(digest_31) : $signed(_GEN_5866); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6370 = 6'h2f == state ? $signed(digest_32) : $signed(_GEN_5867); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6371 = 6'h2f == state ? $signed(digest_33) : $signed(_GEN_5868); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6372 = 6'h2f == state ? $signed(digest_34) : $signed(_GEN_5869); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6373 = 6'h2f == state ? $signed(digest_35) : $signed(_GEN_5870); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6374 = 6'h2f == state ? $signed(digest_36) : $signed(_GEN_5871); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6375 = 6'h2f == state ? $signed(digest_37) : $signed(_GEN_5872); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6376 = 6'h2f == state ? $signed(digest_38) : $signed(_GEN_5873); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6377 = 6'h2f == state ? $signed(digest_39) : $signed(_GEN_5874); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6378 = 6'h2f == state ? $signed(digest_40) : $signed(_GEN_5875); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6379 = 6'h2f == state ? $signed(digest_41) : $signed(_GEN_5876); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6380 = 6'h2f == state ? $signed(digest_42) : $signed(_GEN_5877); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6381 = 6'h2f == state ? $signed(digest_43) : $signed(_GEN_5878); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6382 = 6'h2f == state ? $signed(digest_44) : $signed(_GEN_5879); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6383 = 6'h2f == state ? $signed(digest_45) : $signed(_GEN_5880); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6384 = 6'h2f == state ? $signed(digest_46) : $signed(_GEN_5881); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6385 = 6'h2f == state ? $signed(digest_47) : $signed(_GEN_5882); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6386 = 6'h2f == state ? $signed(digest_48) : $signed(_GEN_5883); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6387 = 6'h2f == state ? $signed(digest_49) : $signed(_GEN_5884); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6388 = 6'h2f == state ? $signed(digest_50) : $signed(_GEN_5885); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6389 = 6'h2f == state ? $signed(digest_51) : $signed(_GEN_5886); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6390 = 6'h2f == state ? $signed(digest_52) : $signed(_GEN_5887); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6391 = 6'h2f == state ? $signed(digest_53) : $signed(_GEN_5888); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6392 = 6'h2f == state ? $signed(digest_54) : $signed(_GEN_5889); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6393 = 6'h2f == state ? $signed(digest_55) : $signed(_GEN_5890); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6394 = 6'h2f == state ? $signed(digest_56) : $signed(_GEN_5891); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6395 = 6'h2f == state ? $signed(digest_57) : $signed(_GEN_5892); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6396 = 6'h2f == state ? $signed(digest_58) : $signed(_GEN_5893); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6397 = 6'h2f == state ? $signed(digest_59) : $signed(_GEN_5894); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6398 = 6'h2f == state ? $signed(digest_60) : $signed(_GEN_5895); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6399 = 6'h2f == state ? $signed(digest_61) : $signed(_GEN_5896); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6400 = 6'h2f == state ? $signed(digest_62) : $signed(_GEN_5897); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6401 = 6'h2f == state ? $signed(digest_63) : $signed(_GEN_5898); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6402 = 6'h2f == state ? $signed(digest_64) : $signed(_GEN_5899); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6403 = 6'h2f == state ? $signed(digest_65) : $signed(_GEN_5900); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6404 = 6'h2f == state ? $signed(digest_66) : $signed(_GEN_5901); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6405 = 6'h2f == state ? $signed(digest_67) : $signed(_GEN_5902); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6406 = 6'h2f == state ? $signed(digest_68) : $signed(_GEN_5903); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6407 = 6'h2f == state ? $signed(digest_69) : $signed(_GEN_5904); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6408 = 6'h2f == state ? $signed(digest_70) : $signed(_GEN_5905); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6409 = 6'h2f == state ? $signed(digest_71) : $signed(_GEN_5906); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6410 = 6'h2f == state ? $signed(digest_72) : $signed(_GEN_5907); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6411 = 6'h2f == state ? $signed(digest_73) : $signed(_GEN_5908); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6412 = 6'h2f == state ? $signed(digest_74) : $signed(_GEN_5909); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6413 = 6'h2f == state ? $signed(digest_75) : $signed(_GEN_5910); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6414 = 6'h2f == state ? $signed(digest_76) : $signed(_GEN_5911); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6415 = 6'h2f == state ? $signed(digest_77) : $signed(_GEN_5912); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6416 = 6'h2f == state ? $signed(digest_78) : $signed(_GEN_5913); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6417 = 6'h2f == state ? $signed(digest_79) : $signed(_GEN_5914); // @[digest.scala 81:19 53:21]
  wire  _GEN_6419 = 6'h2f == state ? 1'h0 : _GEN_5916; // @[digest.scala 81:19 58:25]
  wire  _GEN_6502 = 6'h2f == state ? 1'h0 : _GEN_5999; // @[digest.scala 81:19 63:25]
  wire  _GEN_6585 = 6'h2f == state ? 1'h0 : _GEN_6082; // @[digest.scala 81:19 68:25]
  wire  _GEN_6668 = 6'h2f == state ? 1'h0 : _GEN_6165; // @[digest.scala 81:19 73:25]
  wire  _GEN_6751 = 6'h2f == state ? 1'h0 : _GEN_6248; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_6752 = 6'h2e == state ? $signed(t) : $signed(_GEN_6251); // @[digest.scala 272:15 81:19]
  wire [5:0] _GEN_6753 = 6'h2e == state ? 6'h2f : _GEN_6250; // @[digest.scala 273:19 81:19]
  wire [31:0] _GEN_6754 = 6'h2e == state ? $signed(j) : $signed(_GEN_6249); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_6755 = 6'h2e == state ? $signed(b) : $signed(_GEN_6252); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_6756 = 6'h2e == state ? $signed(c) : $signed(_GEN_6253); // @[digest.scala 26:16 81:19]
  wire [31:0] _GEN_6757 = 6'h2e == state ? $signed(d) : $signed(_GEN_6254); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_6758 = 6'h2e == state ? $signed(e) : $signed(_GEN_6255); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_6759 = 6'h2e == state ? $signed(i) : $signed(_GEN_6256); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_6841 = 6'h2e == state ? $signed(digest_0) : $signed(_GEN_6338); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6842 = 6'h2e == state ? $signed(digest_1) : $signed(_GEN_6339); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6843 = 6'h2e == state ? $signed(digest_2) : $signed(_GEN_6340); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6844 = 6'h2e == state ? $signed(digest_3) : $signed(_GEN_6341); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6845 = 6'h2e == state ? $signed(digest_4) : $signed(_GEN_6342); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6846 = 6'h2e == state ? $signed(digest_5) : $signed(_GEN_6343); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6847 = 6'h2e == state ? $signed(digest_6) : $signed(_GEN_6344); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6848 = 6'h2e == state ? $signed(digest_7) : $signed(_GEN_6345); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6849 = 6'h2e == state ? $signed(digest_8) : $signed(_GEN_6346); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6850 = 6'h2e == state ? $signed(digest_9) : $signed(_GEN_6347); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6851 = 6'h2e == state ? $signed(digest_10) : $signed(_GEN_6348); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6852 = 6'h2e == state ? $signed(digest_11) : $signed(_GEN_6349); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6853 = 6'h2e == state ? $signed(digest_12) : $signed(_GEN_6350); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6854 = 6'h2e == state ? $signed(digest_13) : $signed(_GEN_6351); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6855 = 6'h2e == state ? $signed(digest_14) : $signed(_GEN_6352); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6856 = 6'h2e == state ? $signed(digest_15) : $signed(_GEN_6353); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6857 = 6'h2e == state ? $signed(digest_16) : $signed(_GEN_6354); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6858 = 6'h2e == state ? $signed(digest_17) : $signed(_GEN_6355); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6859 = 6'h2e == state ? $signed(digest_18) : $signed(_GEN_6356); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6860 = 6'h2e == state ? $signed(digest_19) : $signed(_GEN_6357); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6861 = 6'h2e == state ? $signed(digest_20) : $signed(_GEN_6358); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6862 = 6'h2e == state ? $signed(digest_21) : $signed(_GEN_6359); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6863 = 6'h2e == state ? $signed(digest_22) : $signed(_GEN_6360); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6864 = 6'h2e == state ? $signed(digest_23) : $signed(_GEN_6361); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6865 = 6'h2e == state ? $signed(digest_24) : $signed(_GEN_6362); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6866 = 6'h2e == state ? $signed(digest_25) : $signed(_GEN_6363); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6867 = 6'h2e == state ? $signed(digest_26) : $signed(_GEN_6364); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6868 = 6'h2e == state ? $signed(digest_27) : $signed(_GEN_6365); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6869 = 6'h2e == state ? $signed(digest_28) : $signed(_GEN_6366); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6870 = 6'h2e == state ? $signed(digest_29) : $signed(_GEN_6367); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6871 = 6'h2e == state ? $signed(digest_30) : $signed(_GEN_6368); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6872 = 6'h2e == state ? $signed(digest_31) : $signed(_GEN_6369); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6873 = 6'h2e == state ? $signed(digest_32) : $signed(_GEN_6370); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6874 = 6'h2e == state ? $signed(digest_33) : $signed(_GEN_6371); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6875 = 6'h2e == state ? $signed(digest_34) : $signed(_GEN_6372); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6876 = 6'h2e == state ? $signed(digest_35) : $signed(_GEN_6373); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6877 = 6'h2e == state ? $signed(digest_36) : $signed(_GEN_6374); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6878 = 6'h2e == state ? $signed(digest_37) : $signed(_GEN_6375); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6879 = 6'h2e == state ? $signed(digest_38) : $signed(_GEN_6376); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6880 = 6'h2e == state ? $signed(digest_39) : $signed(_GEN_6377); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6881 = 6'h2e == state ? $signed(digest_40) : $signed(_GEN_6378); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6882 = 6'h2e == state ? $signed(digest_41) : $signed(_GEN_6379); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6883 = 6'h2e == state ? $signed(digest_42) : $signed(_GEN_6380); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6884 = 6'h2e == state ? $signed(digest_43) : $signed(_GEN_6381); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6885 = 6'h2e == state ? $signed(digest_44) : $signed(_GEN_6382); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6886 = 6'h2e == state ? $signed(digest_45) : $signed(_GEN_6383); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6887 = 6'h2e == state ? $signed(digest_46) : $signed(_GEN_6384); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6888 = 6'h2e == state ? $signed(digest_47) : $signed(_GEN_6385); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6889 = 6'h2e == state ? $signed(digest_48) : $signed(_GEN_6386); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6890 = 6'h2e == state ? $signed(digest_49) : $signed(_GEN_6387); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6891 = 6'h2e == state ? $signed(digest_50) : $signed(_GEN_6388); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6892 = 6'h2e == state ? $signed(digest_51) : $signed(_GEN_6389); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6893 = 6'h2e == state ? $signed(digest_52) : $signed(_GEN_6390); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6894 = 6'h2e == state ? $signed(digest_53) : $signed(_GEN_6391); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6895 = 6'h2e == state ? $signed(digest_54) : $signed(_GEN_6392); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6896 = 6'h2e == state ? $signed(digest_55) : $signed(_GEN_6393); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6897 = 6'h2e == state ? $signed(digest_56) : $signed(_GEN_6394); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6898 = 6'h2e == state ? $signed(digest_57) : $signed(_GEN_6395); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6899 = 6'h2e == state ? $signed(digest_58) : $signed(_GEN_6396); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6900 = 6'h2e == state ? $signed(digest_59) : $signed(_GEN_6397); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6901 = 6'h2e == state ? $signed(digest_60) : $signed(_GEN_6398); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6902 = 6'h2e == state ? $signed(digest_61) : $signed(_GEN_6399); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6903 = 6'h2e == state ? $signed(digest_62) : $signed(_GEN_6400); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6904 = 6'h2e == state ? $signed(digest_63) : $signed(_GEN_6401); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6905 = 6'h2e == state ? $signed(digest_64) : $signed(_GEN_6402); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6906 = 6'h2e == state ? $signed(digest_65) : $signed(_GEN_6403); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6907 = 6'h2e == state ? $signed(digest_66) : $signed(_GEN_6404); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6908 = 6'h2e == state ? $signed(digest_67) : $signed(_GEN_6405); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6909 = 6'h2e == state ? $signed(digest_68) : $signed(_GEN_6406); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6910 = 6'h2e == state ? $signed(digest_69) : $signed(_GEN_6407); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6911 = 6'h2e == state ? $signed(digest_70) : $signed(_GEN_6408); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6912 = 6'h2e == state ? $signed(digest_71) : $signed(_GEN_6409); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6913 = 6'h2e == state ? $signed(digest_72) : $signed(_GEN_6410); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6914 = 6'h2e == state ? $signed(digest_73) : $signed(_GEN_6411); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6915 = 6'h2e == state ? $signed(digest_74) : $signed(_GEN_6412); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6916 = 6'h2e == state ? $signed(digest_75) : $signed(_GEN_6413); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6917 = 6'h2e == state ? $signed(digest_76) : $signed(_GEN_6414); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6918 = 6'h2e == state ? $signed(digest_77) : $signed(_GEN_6415); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6919 = 6'h2e == state ? $signed(digest_78) : $signed(_GEN_6416); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_6920 = 6'h2e == state ? $signed(digest_79) : $signed(_GEN_6417); // @[digest.scala 81:19 53:21]
  wire  _GEN_6922 = 6'h2e == state ? 1'h0 : _GEN_6419; // @[digest.scala 81:19 58:25]
  wire  _GEN_7005 = 6'h2e == state ? 1'h0 : _GEN_6502; // @[digest.scala 81:19 63:25]
  wire  _GEN_7088 = 6'h2e == state ? 1'h0 : _GEN_6585; // @[digest.scala 81:19 68:25]
  wire  _GEN_7171 = 6'h2e == state ? 1'h0 : _GEN_6668; // @[digest.scala 81:19 73:25]
  wire  _GEN_7254 = 6'h2e == state ? 1'h0 : _GEN_6751; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_7255 = 6'h2d == state ? $signed(a) : $signed(_GEN_6755); // @[digest.scala 268:15 81:19]
  wire [5:0] _GEN_7256 = 6'h2d == state ? 6'h2e : _GEN_6753; // @[digest.scala 269:19 81:19]
  wire [31:0] _GEN_7257 = 6'h2d == state ? $signed(a) : $signed(_GEN_6752); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_7258 = 6'h2d == state ? $signed(j) : $signed(_GEN_6754); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_7259 = 6'h2d == state ? $signed(c) : $signed(_GEN_6756); // @[digest.scala 26:16 81:19]
  wire [31:0] _GEN_7260 = 6'h2d == state ? $signed(d) : $signed(_GEN_6757); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_7261 = 6'h2d == state ? $signed(e) : $signed(_GEN_6758); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_7262 = 6'h2d == state ? $signed(i) : $signed(_GEN_6759); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_7344 = 6'h2d == state ? $signed(digest_0) : $signed(_GEN_6841); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7345 = 6'h2d == state ? $signed(digest_1) : $signed(_GEN_6842); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7346 = 6'h2d == state ? $signed(digest_2) : $signed(_GEN_6843); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7347 = 6'h2d == state ? $signed(digest_3) : $signed(_GEN_6844); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7348 = 6'h2d == state ? $signed(digest_4) : $signed(_GEN_6845); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7349 = 6'h2d == state ? $signed(digest_5) : $signed(_GEN_6846); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7350 = 6'h2d == state ? $signed(digest_6) : $signed(_GEN_6847); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7351 = 6'h2d == state ? $signed(digest_7) : $signed(_GEN_6848); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7352 = 6'h2d == state ? $signed(digest_8) : $signed(_GEN_6849); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7353 = 6'h2d == state ? $signed(digest_9) : $signed(_GEN_6850); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7354 = 6'h2d == state ? $signed(digest_10) : $signed(_GEN_6851); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7355 = 6'h2d == state ? $signed(digest_11) : $signed(_GEN_6852); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7356 = 6'h2d == state ? $signed(digest_12) : $signed(_GEN_6853); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7357 = 6'h2d == state ? $signed(digest_13) : $signed(_GEN_6854); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7358 = 6'h2d == state ? $signed(digest_14) : $signed(_GEN_6855); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7359 = 6'h2d == state ? $signed(digest_15) : $signed(_GEN_6856); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7360 = 6'h2d == state ? $signed(digest_16) : $signed(_GEN_6857); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7361 = 6'h2d == state ? $signed(digest_17) : $signed(_GEN_6858); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7362 = 6'h2d == state ? $signed(digest_18) : $signed(_GEN_6859); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7363 = 6'h2d == state ? $signed(digest_19) : $signed(_GEN_6860); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7364 = 6'h2d == state ? $signed(digest_20) : $signed(_GEN_6861); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7365 = 6'h2d == state ? $signed(digest_21) : $signed(_GEN_6862); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7366 = 6'h2d == state ? $signed(digest_22) : $signed(_GEN_6863); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7367 = 6'h2d == state ? $signed(digest_23) : $signed(_GEN_6864); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7368 = 6'h2d == state ? $signed(digest_24) : $signed(_GEN_6865); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7369 = 6'h2d == state ? $signed(digest_25) : $signed(_GEN_6866); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7370 = 6'h2d == state ? $signed(digest_26) : $signed(_GEN_6867); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7371 = 6'h2d == state ? $signed(digest_27) : $signed(_GEN_6868); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7372 = 6'h2d == state ? $signed(digest_28) : $signed(_GEN_6869); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7373 = 6'h2d == state ? $signed(digest_29) : $signed(_GEN_6870); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7374 = 6'h2d == state ? $signed(digest_30) : $signed(_GEN_6871); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7375 = 6'h2d == state ? $signed(digest_31) : $signed(_GEN_6872); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7376 = 6'h2d == state ? $signed(digest_32) : $signed(_GEN_6873); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7377 = 6'h2d == state ? $signed(digest_33) : $signed(_GEN_6874); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7378 = 6'h2d == state ? $signed(digest_34) : $signed(_GEN_6875); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7379 = 6'h2d == state ? $signed(digest_35) : $signed(_GEN_6876); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7380 = 6'h2d == state ? $signed(digest_36) : $signed(_GEN_6877); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7381 = 6'h2d == state ? $signed(digest_37) : $signed(_GEN_6878); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7382 = 6'h2d == state ? $signed(digest_38) : $signed(_GEN_6879); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7383 = 6'h2d == state ? $signed(digest_39) : $signed(_GEN_6880); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7384 = 6'h2d == state ? $signed(digest_40) : $signed(_GEN_6881); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7385 = 6'h2d == state ? $signed(digest_41) : $signed(_GEN_6882); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7386 = 6'h2d == state ? $signed(digest_42) : $signed(_GEN_6883); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7387 = 6'h2d == state ? $signed(digest_43) : $signed(_GEN_6884); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7388 = 6'h2d == state ? $signed(digest_44) : $signed(_GEN_6885); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7389 = 6'h2d == state ? $signed(digest_45) : $signed(_GEN_6886); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7390 = 6'h2d == state ? $signed(digest_46) : $signed(_GEN_6887); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7391 = 6'h2d == state ? $signed(digest_47) : $signed(_GEN_6888); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7392 = 6'h2d == state ? $signed(digest_48) : $signed(_GEN_6889); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7393 = 6'h2d == state ? $signed(digest_49) : $signed(_GEN_6890); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7394 = 6'h2d == state ? $signed(digest_50) : $signed(_GEN_6891); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7395 = 6'h2d == state ? $signed(digest_51) : $signed(_GEN_6892); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7396 = 6'h2d == state ? $signed(digest_52) : $signed(_GEN_6893); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7397 = 6'h2d == state ? $signed(digest_53) : $signed(_GEN_6894); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7398 = 6'h2d == state ? $signed(digest_54) : $signed(_GEN_6895); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7399 = 6'h2d == state ? $signed(digest_55) : $signed(_GEN_6896); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7400 = 6'h2d == state ? $signed(digest_56) : $signed(_GEN_6897); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7401 = 6'h2d == state ? $signed(digest_57) : $signed(_GEN_6898); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7402 = 6'h2d == state ? $signed(digest_58) : $signed(_GEN_6899); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7403 = 6'h2d == state ? $signed(digest_59) : $signed(_GEN_6900); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7404 = 6'h2d == state ? $signed(digest_60) : $signed(_GEN_6901); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7405 = 6'h2d == state ? $signed(digest_61) : $signed(_GEN_6902); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7406 = 6'h2d == state ? $signed(digest_62) : $signed(_GEN_6903); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7407 = 6'h2d == state ? $signed(digest_63) : $signed(_GEN_6904); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7408 = 6'h2d == state ? $signed(digest_64) : $signed(_GEN_6905); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7409 = 6'h2d == state ? $signed(digest_65) : $signed(_GEN_6906); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7410 = 6'h2d == state ? $signed(digest_66) : $signed(_GEN_6907); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7411 = 6'h2d == state ? $signed(digest_67) : $signed(_GEN_6908); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7412 = 6'h2d == state ? $signed(digest_68) : $signed(_GEN_6909); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7413 = 6'h2d == state ? $signed(digest_69) : $signed(_GEN_6910); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7414 = 6'h2d == state ? $signed(digest_70) : $signed(_GEN_6911); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7415 = 6'h2d == state ? $signed(digest_71) : $signed(_GEN_6912); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7416 = 6'h2d == state ? $signed(digest_72) : $signed(_GEN_6913); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7417 = 6'h2d == state ? $signed(digest_73) : $signed(_GEN_6914); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7418 = 6'h2d == state ? $signed(digest_74) : $signed(_GEN_6915); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7419 = 6'h2d == state ? $signed(digest_75) : $signed(_GEN_6916); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7420 = 6'h2d == state ? $signed(digest_76) : $signed(_GEN_6917); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7421 = 6'h2d == state ? $signed(digest_77) : $signed(_GEN_6918); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7422 = 6'h2d == state ? $signed(digest_78) : $signed(_GEN_6919); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7423 = 6'h2d == state ? $signed(digest_79) : $signed(_GEN_6920); // @[digest.scala 81:19 53:21]
  wire  _GEN_7425 = 6'h2d == state ? 1'h0 : _GEN_6922; // @[digest.scala 81:19 58:25]
  wire  _GEN_7508 = 6'h2d == state ? 1'h0 : _GEN_7005; // @[digest.scala 81:19 63:25]
  wire  _GEN_7591 = 6'h2d == state ? 1'h0 : _GEN_7088; // @[digest.scala 81:19 68:25]
  wire  _GEN_7674 = 6'h2d == state ? 1'h0 : _GEN_7171; // @[digest.scala 81:19 73:25]
  wire  _GEN_7757 = 6'h2d == state ? 1'h0 : _GEN_7254; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_7758 = 6'h2c == state ? $signed(__m_rol_2_io_out_rol) : $signed(_GEN_7259); // @[digest.scala 261:15 81:19]
  wire  _GEN_7759 = 6'h2c == state & __m_rol_2_io_valid_T; // @[digest.scala 81:19 262:32 52:24]
  wire [5:0] _GEN_7762 = 6'h2c == state ? _state_T_17 : _GEN_7256; // @[digest.scala 265:19 81:19]
  wire [31:0] _GEN_7763 = 6'h2c == state ? $signed(b) : $signed(_GEN_7255); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_7764 = 6'h2c == state ? $signed(a) : $signed(_GEN_7257); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_7765 = 6'h2c == state ? $signed(j) : $signed(_GEN_7258); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_7766 = 6'h2c == state ? $signed(d) : $signed(_GEN_7260); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_7767 = 6'h2c == state ? $signed(e) : $signed(_GEN_7261); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_7768 = 6'h2c == state ? $signed(i) : $signed(_GEN_7262); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_7850 = 6'h2c == state ? $signed(digest_0) : $signed(_GEN_7344); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7851 = 6'h2c == state ? $signed(digest_1) : $signed(_GEN_7345); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7852 = 6'h2c == state ? $signed(digest_2) : $signed(_GEN_7346); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7853 = 6'h2c == state ? $signed(digest_3) : $signed(_GEN_7347); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7854 = 6'h2c == state ? $signed(digest_4) : $signed(_GEN_7348); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7855 = 6'h2c == state ? $signed(digest_5) : $signed(_GEN_7349); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7856 = 6'h2c == state ? $signed(digest_6) : $signed(_GEN_7350); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7857 = 6'h2c == state ? $signed(digest_7) : $signed(_GEN_7351); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7858 = 6'h2c == state ? $signed(digest_8) : $signed(_GEN_7352); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7859 = 6'h2c == state ? $signed(digest_9) : $signed(_GEN_7353); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7860 = 6'h2c == state ? $signed(digest_10) : $signed(_GEN_7354); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7861 = 6'h2c == state ? $signed(digest_11) : $signed(_GEN_7355); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7862 = 6'h2c == state ? $signed(digest_12) : $signed(_GEN_7356); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7863 = 6'h2c == state ? $signed(digest_13) : $signed(_GEN_7357); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7864 = 6'h2c == state ? $signed(digest_14) : $signed(_GEN_7358); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7865 = 6'h2c == state ? $signed(digest_15) : $signed(_GEN_7359); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7866 = 6'h2c == state ? $signed(digest_16) : $signed(_GEN_7360); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7867 = 6'h2c == state ? $signed(digest_17) : $signed(_GEN_7361); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7868 = 6'h2c == state ? $signed(digest_18) : $signed(_GEN_7362); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7869 = 6'h2c == state ? $signed(digest_19) : $signed(_GEN_7363); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7870 = 6'h2c == state ? $signed(digest_20) : $signed(_GEN_7364); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7871 = 6'h2c == state ? $signed(digest_21) : $signed(_GEN_7365); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7872 = 6'h2c == state ? $signed(digest_22) : $signed(_GEN_7366); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7873 = 6'h2c == state ? $signed(digest_23) : $signed(_GEN_7367); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7874 = 6'h2c == state ? $signed(digest_24) : $signed(_GEN_7368); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7875 = 6'h2c == state ? $signed(digest_25) : $signed(_GEN_7369); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7876 = 6'h2c == state ? $signed(digest_26) : $signed(_GEN_7370); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7877 = 6'h2c == state ? $signed(digest_27) : $signed(_GEN_7371); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7878 = 6'h2c == state ? $signed(digest_28) : $signed(_GEN_7372); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7879 = 6'h2c == state ? $signed(digest_29) : $signed(_GEN_7373); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7880 = 6'h2c == state ? $signed(digest_30) : $signed(_GEN_7374); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7881 = 6'h2c == state ? $signed(digest_31) : $signed(_GEN_7375); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7882 = 6'h2c == state ? $signed(digest_32) : $signed(_GEN_7376); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7883 = 6'h2c == state ? $signed(digest_33) : $signed(_GEN_7377); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7884 = 6'h2c == state ? $signed(digest_34) : $signed(_GEN_7378); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7885 = 6'h2c == state ? $signed(digest_35) : $signed(_GEN_7379); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7886 = 6'h2c == state ? $signed(digest_36) : $signed(_GEN_7380); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7887 = 6'h2c == state ? $signed(digest_37) : $signed(_GEN_7381); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7888 = 6'h2c == state ? $signed(digest_38) : $signed(_GEN_7382); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7889 = 6'h2c == state ? $signed(digest_39) : $signed(_GEN_7383); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7890 = 6'h2c == state ? $signed(digest_40) : $signed(_GEN_7384); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7891 = 6'h2c == state ? $signed(digest_41) : $signed(_GEN_7385); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7892 = 6'h2c == state ? $signed(digest_42) : $signed(_GEN_7386); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7893 = 6'h2c == state ? $signed(digest_43) : $signed(_GEN_7387); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7894 = 6'h2c == state ? $signed(digest_44) : $signed(_GEN_7388); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7895 = 6'h2c == state ? $signed(digest_45) : $signed(_GEN_7389); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7896 = 6'h2c == state ? $signed(digest_46) : $signed(_GEN_7390); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7897 = 6'h2c == state ? $signed(digest_47) : $signed(_GEN_7391); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7898 = 6'h2c == state ? $signed(digest_48) : $signed(_GEN_7392); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7899 = 6'h2c == state ? $signed(digest_49) : $signed(_GEN_7393); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7900 = 6'h2c == state ? $signed(digest_50) : $signed(_GEN_7394); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7901 = 6'h2c == state ? $signed(digest_51) : $signed(_GEN_7395); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7902 = 6'h2c == state ? $signed(digest_52) : $signed(_GEN_7396); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7903 = 6'h2c == state ? $signed(digest_53) : $signed(_GEN_7397); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7904 = 6'h2c == state ? $signed(digest_54) : $signed(_GEN_7398); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7905 = 6'h2c == state ? $signed(digest_55) : $signed(_GEN_7399); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7906 = 6'h2c == state ? $signed(digest_56) : $signed(_GEN_7400); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7907 = 6'h2c == state ? $signed(digest_57) : $signed(_GEN_7401); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7908 = 6'h2c == state ? $signed(digest_58) : $signed(_GEN_7402); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7909 = 6'h2c == state ? $signed(digest_59) : $signed(_GEN_7403); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7910 = 6'h2c == state ? $signed(digest_60) : $signed(_GEN_7404); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7911 = 6'h2c == state ? $signed(digest_61) : $signed(_GEN_7405); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7912 = 6'h2c == state ? $signed(digest_62) : $signed(_GEN_7406); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7913 = 6'h2c == state ? $signed(digest_63) : $signed(_GEN_7407); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7914 = 6'h2c == state ? $signed(digest_64) : $signed(_GEN_7408); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7915 = 6'h2c == state ? $signed(digest_65) : $signed(_GEN_7409); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7916 = 6'h2c == state ? $signed(digest_66) : $signed(_GEN_7410); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7917 = 6'h2c == state ? $signed(digest_67) : $signed(_GEN_7411); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7918 = 6'h2c == state ? $signed(digest_68) : $signed(_GEN_7412); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7919 = 6'h2c == state ? $signed(digest_69) : $signed(_GEN_7413); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7920 = 6'h2c == state ? $signed(digest_70) : $signed(_GEN_7414); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7921 = 6'h2c == state ? $signed(digest_71) : $signed(_GEN_7415); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7922 = 6'h2c == state ? $signed(digest_72) : $signed(_GEN_7416); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7923 = 6'h2c == state ? $signed(digest_73) : $signed(_GEN_7417); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7924 = 6'h2c == state ? $signed(digest_74) : $signed(_GEN_7418); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7925 = 6'h2c == state ? $signed(digest_75) : $signed(_GEN_7419); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7926 = 6'h2c == state ? $signed(digest_76) : $signed(_GEN_7420); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7927 = 6'h2c == state ? $signed(digest_77) : $signed(_GEN_7421); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7928 = 6'h2c == state ? $signed(digest_78) : $signed(_GEN_7422); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_7929 = 6'h2c == state ? $signed(digest_79) : $signed(_GEN_7423); // @[digest.scala 81:19 53:21]
  wire  _GEN_7931 = 6'h2c == state ? 1'h0 : _GEN_7425; // @[digest.scala 81:19 58:25]
  wire  _GEN_8014 = 6'h2c == state ? 1'h0 : _GEN_7508; // @[digest.scala 81:19 63:25]
  wire  _GEN_8097 = 6'h2c == state ? 1'h0 : _GEN_7591; // @[digest.scala 81:19 68:25]
  wire  _GEN_8180 = 6'h2c == state ? 1'h0 : _GEN_7674; // @[digest.scala 81:19 73:25]
  wire  _GEN_8263 = 6'h2c == state ? 1'h0 : _GEN_7757; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_8264 = 6'h2b == state ? $signed(c) : $signed(_GEN_7766); // @[digest.scala 257:15 81:19]
  wire [5:0] _GEN_8265 = 6'h2b == state ? 6'h2c : _GEN_7762; // @[digest.scala 258:19 81:19]
  wire [31:0] _GEN_8266 = 6'h2b == state ? $signed(c) : $signed(_GEN_7758); // @[digest.scala 26:16 81:19]
  wire  _GEN_8267 = 6'h2b == state ? 1'h0 : _GEN_7759; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_8270 = 6'h2b == state ? $signed(b) : $signed(_GEN_7763); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_8271 = 6'h2b == state ? $signed(a) : $signed(_GEN_7764); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_8272 = 6'h2b == state ? $signed(j) : $signed(_GEN_7765); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_8273 = 6'h2b == state ? $signed(e) : $signed(_GEN_7767); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_8274 = 6'h2b == state ? $signed(i) : $signed(_GEN_7768); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_8356 = 6'h2b == state ? $signed(digest_0) : $signed(_GEN_7850); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8357 = 6'h2b == state ? $signed(digest_1) : $signed(_GEN_7851); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8358 = 6'h2b == state ? $signed(digest_2) : $signed(_GEN_7852); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8359 = 6'h2b == state ? $signed(digest_3) : $signed(_GEN_7853); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8360 = 6'h2b == state ? $signed(digest_4) : $signed(_GEN_7854); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8361 = 6'h2b == state ? $signed(digest_5) : $signed(_GEN_7855); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8362 = 6'h2b == state ? $signed(digest_6) : $signed(_GEN_7856); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8363 = 6'h2b == state ? $signed(digest_7) : $signed(_GEN_7857); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8364 = 6'h2b == state ? $signed(digest_8) : $signed(_GEN_7858); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8365 = 6'h2b == state ? $signed(digest_9) : $signed(_GEN_7859); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8366 = 6'h2b == state ? $signed(digest_10) : $signed(_GEN_7860); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8367 = 6'h2b == state ? $signed(digest_11) : $signed(_GEN_7861); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8368 = 6'h2b == state ? $signed(digest_12) : $signed(_GEN_7862); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8369 = 6'h2b == state ? $signed(digest_13) : $signed(_GEN_7863); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8370 = 6'h2b == state ? $signed(digest_14) : $signed(_GEN_7864); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8371 = 6'h2b == state ? $signed(digest_15) : $signed(_GEN_7865); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8372 = 6'h2b == state ? $signed(digest_16) : $signed(_GEN_7866); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8373 = 6'h2b == state ? $signed(digest_17) : $signed(_GEN_7867); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8374 = 6'h2b == state ? $signed(digest_18) : $signed(_GEN_7868); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8375 = 6'h2b == state ? $signed(digest_19) : $signed(_GEN_7869); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8376 = 6'h2b == state ? $signed(digest_20) : $signed(_GEN_7870); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8377 = 6'h2b == state ? $signed(digest_21) : $signed(_GEN_7871); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8378 = 6'h2b == state ? $signed(digest_22) : $signed(_GEN_7872); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8379 = 6'h2b == state ? $signed(digest_23) : $signed(_GEN_7873); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8380 = 6'h2b == state ? $signed(digest_24) : $signed(_GEN_7874); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8381 = 6'h2b == state ? $signed(digest_25) : $signed(_GEN_7875); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8382 = 6'h2b == state ? $signed(digest_26) : $signed(_GEN_7876); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8383 = 6'h2b == state ? $signed(digest_27) : $signed(_GEN_7877); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8384 = 6'h2b == state ? $signed(digest_28) : $signed(_GEN_7878); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8385 = 6'h2b == state ? $signed(digest_29) : $signed(_GEN_7879); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8386 = 6'h2b == state ? $signed(digest_30) : $signed(_GEN_7880); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8387 = 6'h2b == state ? $signed(digest_31) : $signed(_GEN_7881); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8388 = 6'h2b == state ? $signed(digest_32) : $signed(_GEN_7882); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8389 = 6'h2b == state ? $signed(digest_33) : $signed(_GEN_7883); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8390 = 6'h2b == state ? $signed(digest_34) : $signed(_GEN_7884); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8391 = 6'h2b == state ? $signed(digest_35) : $signed(_GEN_7885); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8392 = 6'h2b == state ? $signed(digest_36) : $signed(_GEN_7886); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8393 = 6'h2b == state ? $signed(digest_37) : $signed(_GEN_7887); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8394 = 6'h2b == state ? $signed(digest_38) : $signed(_GEN_7888); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8395 = 6'h2b == state ? $signed(digest_39) : $signed(_GEN_7889); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8396 = 6'h2b == state ? $signed(digest_40) : $signed(_GEN_7890); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8397 = 6'h2b == state ? $signed(digest_41) : $signed(_GEN_7891); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8398 = 6'h2b == state ? $signed(digest_42) : $signed(_GEN_7892); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8399 = 6'h2b == state ? $signed(digest_43) : $signed(_GEN_7893); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8400 = 6'h2b == state ? $signed(digest_44) : $signed(_GEN_7894); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8401 = 6'h2b == state ? $signed(digest_45) : $signed(_GEN_7895); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8402 = 6'h2b == state ? $signed(digest_46) : $signed(_GEN_7896); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8403 = 6'h2b == state ? $signed(digest_47) : $signed(_GEN_7897); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8404 = 6'h2b == state ? $signed(digest_48) : $signed(_GEN_7898); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8405 = 6'h2b == state ? $signed(digest_49) : $signed(_GEN_7899); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8406 = 6'h2b == state ? $signed(digest_50) : $signed(_GEN_7900); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8407 = 6'h2b == state ? $signed(digest_51) : $signed(_GEN_7901); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8408 = 6'h2b == state ? $signed(digest_52) : $signed(_GEN_7902); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8409 = 6'h2b == state ? $signed(digest_53) : $signed(_GEN_7903); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8410 = 6'h2b == state ? $signed(digest_54) : $signed(_GEN_7904); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8411 = 6'h2b == state ? $signed(digest_55) : $signed(_GEN_7905); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8412 = 6'h2b == state ? $signed(digest_56) : $signed(_GEN_7906); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8413 = 6'h2b == state ? $signed(digest_57) : $signed(_GEN_7907); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8414 = 6'h2b == state ? $signed(digest_58) : $signed(_GEN_7908); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8415 = 6'h2b == state ? $signed(digest_59) : $signed(_GEN_7909); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8416 = 6'h2b == state ? $signed(digest_60) : $signed(_GEN_7910); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8417 = 6'h2b == state ? $signed(digest_61) : $signed(_GEN_7911); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8418 = 6'h2b == state ? $signed(digest_62) : $signed(_GEN_7912); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8419 = 6'h2b == state ? $signed(digest_63) : $signed(_GEN_7913); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8420 = 6'h2b == state ? $signed(digest_64) : $signed(_GEN_7914); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8421 = 6'h2b == state ? $signed(digest_65) : $signed(_GEN_7915); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8422 = 6'h2b == state ? $signed(digest_66) : $signed(_GEN_7916); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8423 = 6'h2b == state ? $signed(digest_67) : $signed(_GEN_7917); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8424 = 6'h2b == state ? $signed(digest_68) : $signed(_GEN_7918); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8425 = 6'h2b == state ? $signed(digest_69) : $signed(_GEN_7919); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8426 = 6'h2b == state ? $signed(digest_70) : $signed(_GEN_7920); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8427 = 6'h2b == state ? $signed(digest_71) : $signed(_GEN_7921); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8428 = 6'h2b == state ? $signed(digest_72) : $signed(_GEN_7922); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8429 = 6'h2b == state ? $signed(digest_73) : $signed(_GEN_7923); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8430 = 6'h2b == state ? $signed(digest_74) : $signed(_GEN_7924); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8431 = 6'h2b == state ? $signed(digest_75) : $signed(_GEN_7925); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8432 = 6'h2b == state ? $signed(digest_76) : $signed(_GEN_7926); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8433 = 6'h2b == state ? $signed(digest_77) : $signed(_GEN_7927); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8434 = 6'h2b == state ? $signed(digest_78) : $signed(_GEN_7928); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8435 = 6'h2b == state ? $signed(digest_79) : $signed(_GEN_7929); // @[digest.scala 81:19 53:21]
  wire  _GEN_8437 = 6'h2b == state ? 1'h0 : _GEN_7931; // @[digest.scala 81:19 58:25]
  wire  _GEN_8520 = 6'h2b == state ? 1'h0 : _GEN_8014; // @[digest.scala 81:19 63:25]
  wire  _GEN_8603 = 6'h2b == state ? 1'h0 : _GEN_8097; // @[digest.scala 81:19 68:25]
  wire  _GEN_8686 = 6'h2b == state ? 1'h0 : _GEN_8180; // @[digest.scala 81:19 73:25]
  wire  _GEN_8769 = 6'h2b == state ? 1'h0 : _GEN_8263; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_8770 = 6'h2a == state ? $signed(d) : $signed(_GEN_8273); // @[digest.scala 253:15 81:19]
  wire [5:0] _GEN_8771 = 6'h2a == state ? 6'h2b : _GEN_8265; // @[digest.scala 254:19 81:19]
  wire [31:0] _GEN_8772 = 6'h2a == state ? $signed(d) : $signed(_GEN_8264); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_8773 = 6'h2a == state ? $signed(c) : $signed(_GEN_8266); // @[digest.scala 26:16 81:19]
  wire  _GEN_8774 = 6'h2a == state ? 1'h0 : _GEN_8267; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_8777 = 6'h2a == state ? $signed(b) : $signed(_GEN_8270); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_8778 = 6'h2a == state ? $signed(a) : $signed(_GEN_8271); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_8779 = 6'h2a == state ? $signed(j) : $signed(_GEN_8272); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_8780 = 6'h2a == state ? $signed(i) : $signed(_GEN_8274); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_8862 = 6'h2a == state ? $signed(digest_0) : $signed(_GEN_8356); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8863 = 6'h2a == state ? $signed(digest_1) : $signed(_GEN_8357); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8864 = 6'h2a == state ? $signed(digest_2) : $signed(_GEN_8358); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8865 = 6'h2a == state ? $signed(digest_3) : $signed(_GEN_8359); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8866 = 6'h2a == state ? $signed(digest_4) : $signed(_GEN_8360); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8867 = 6'h2a == state ? $signed(digest_5) : $signed(_GEN_8361); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8868 = 6'h2a == state ? $signed(digest_6) : $signed(_GEN_8362); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8869 = 6'h2a == state ? $signed(digest_7) : $signed(_GEN_8363); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8870 = 6'h2a == state ? $signed(digest_8) : $signed(_GEN_8364); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8871 = 6'h2a == state ? $signed(digest_9) : $signed(_GEN_8365); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8872 = 6'h2a == state ? $signed(digest_10) : $signed(_GEN_8366); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8873 = 6'h2a == state ? $signed(digest_11) : $signed(_GEN_8367); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8874 = 6'h2a == state ? $signed(digest_12) : $signed(_GEN_8368); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8875 = 6'h2a == state ? $signed(digest_13) : $signed(_GEN_8369); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8876 = 6'h2a == state ? $signed(digest_14) : $signed(_GEN_8370); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8877 = 6'h2a == state ? $signed(digest_15) : $signed(_GEN_8371); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8878 = 6'h2a == state ? $signed(digest_16) : $signed(_GEN_8372); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8879 = 6'h2a == state ? $signed(digest_17) : $signed(_GEN_8373); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8880 = 6'h2a == state ? $signed(digest_18) : $signed(_GEN_8374); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8881 = 6'h2a == state ? $signed(digest_19) : $signed(_GEN_8375); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8882 = 6'h2a == state ? $signed(digest_20) : $signed(_GEN_8376); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8883 = 6'h2a == state ? $signed(digest_21) : $signed(_GEN_8377); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8884 = 6'h2a == state ? $signed(digest_22) : $signed(_GEN_8378); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8885 = 6'h2a == state ? $signed(digest_23) : $signed(_GEN_8379); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8886 = 6'h2a == state ? $signed(digest_24) : $signed(_GEN_8380); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8887 = 6'h2a == state ? $signed(digest_25) : $signed(_GEN_8381); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8888 = 6'h2a == state ? $signed(digest_26) : $signed(_GEN_8382); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8889 = 6'h2a == state ? $signed(digest_27) : $signed(_GEN_8383); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8890 = 6'h2a == state ? $signed(digest_28) : $signed(_GEN_8384); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8891 = 6'h2a == state ? $signed(digest_29) : $signed(_GEN_8385); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8892 = 6'h2a == state ? $signed(digest_30) : $signed(_GEN_8386); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8893 = 6'h2a == state ? $signed(digest_31) : $signed(_GEN_8387); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8894 = 6'h2a == state ? $signed(digest_32) : $signed(_GEN_8388); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8895 = 6'h2a == state ? $signed(digest_33) : $signed(_GEN_8389); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8896 = 6'h2a == state ? $signed(digest_34) : $signed(_GEN_8390); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8897 = 6'h2a == state ? $signed(digest_35) : $signed(_GEN_8391); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8898 = 6'h2a == state ? $signed(digest_36) : $signed(_GEN_8392); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8899 = 6'h2a == state ? $signed(digest_37) : $signed(_GEN_8393); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8900 = 6'h2a == state ? $signed(digest_38) : $signed(_GEN_8394); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8901 = 6'h2a == state ? $signed(digest_39) : $signed(_GEN_8395); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8902 = 6'h2a == state ? $signed(digest_40) : $signed(_GEN_8396); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8903 = 6'h2a == state ? $signed(digest_41) : $signed(_GEN_8397); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8904 = 6'h2a == state ? $signed(digest_42) : $signed(_GEN_8398); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8905 = 6'h2a == state ? $signed(digest_43) : $signed(_GEN_8399); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8906 = 6'h2a == state ? $signed(digest_44) : $signed(_GEN_8400); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8907 = 6'h2a == state ? $signed(digest_45) : $signed(_GEN_8401); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8908 = 6'h2a == state ? $signed(digest_46) : $signed(_GEN_8402); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8909 = 6'h2a == state ? $signed(digest_47) : $signed(_GEN_8403); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8910 = 6'h2a == state ? $signed(digest_48) : $signed(_GEN_8404); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8911 = 6'h2a == state ? $signed(digest_49) : $signed(_GEN_8405); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8912 = 6'h2a == state ? $signed(digest_50) : $signed(_GEN_8406); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8913 = 6'h2a == state ? $signed(digest_51) : $signed(_GEN_8407); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8914 = 6'h2a == state ? $signed(digest_52) : $signed(_GEN_8408); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8915 = 6'h2a == state ? $signed(digest_53) : $signed(_GEN_8409); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8916 = 6'h2a == state ? $signed(digest_54) : $signed(_GEN_8410); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8917 = 6'h2a == state ? $signed(digest_55) : $signed(_GEN_8411); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8918 = 6'h2a == state ? $signed(digest_56) : $signed(_GEN_8412); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8919 = 6'h2a == state ? $signed(digest_57) : $signed(_GEN_8413); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8920 = 6'h2a == state ? $signed(digest_58) : $signed(_GEN_8414); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8921 = 6'h2a == state ? $signed(digest_59) : $signed(_GEN_8415); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8922 = 6'h2a == state ? $signed(digest_60) : $signed(_GEN_8416); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8923 = 6'h2a == state ? $signed(digest_61) : $signed(_GEN_8417); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8924 = 6'h2a == state ? $signed(digest_62) : $signed(_GEN_8418); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8925 = 6'h2a == state ? $signed(digest_63) : $signed(_GEN_8419); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8926 = 6'h2a == state ? $signed(digest_64) : $signed(_GEN_8420); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8927 = 6'h2a == state ? $signed(digest_65) : $signed(_GEN_8421); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8928 = 6'h2a == state ? $signed(digest_66) : $signed(_GEN_8422); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8929 = 6'h2a == state ? $signed(digest_67) : $signed(_GEN_8423); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8930 = 6'h2a == state ? $signed(digest_68) : $signed(_GEN_8424); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8931 = 6'h2a == state ? $signed(digest_69) : $signed(_GEN_8425); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8932 = 6'h2a == state ? $signed(digest_70) : $signed(_GEN_8426); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8933 = 6'h2a == state ? $signed(digest_71) : $signed(_GEN_8427); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8934 = 6'h2a == state ? $signed(digest_72) : $signed(_GEN_8428); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8935 = 6'h2a == state ? $signed(digest_73) : $signed(_GEN_8429); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8936 = 6'h2a == state ? $signed(digest_74) : $signed(_GEN_8430); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8937 = 6'h2a == state ? $signed(digest_75) : $signed(_GEN_8431); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8938 = 6'h2a == state ? $signed(digest_76) : $signed(_GEN_8432); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8939 = 6'h2a == state ? $signed(digest_77) : $signed(_GEN_8433); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8940 = 6'h2a == state ? $signed(digest_78) : $signed(_GEN_8434); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_8941 = 6'h2a == state ? $signed(digest_79) : $signed(_GEN_8435); // @[digest.scala 81:19 53:21]
  wire  _GEN_8943 = 6'h2a == state ? 1'h0 : _GEN_8437; // @[digest.scala 81:19 58:25]
  wire  _GEN_9026 = 6'h2a == state ? 1'h0 : _GEN_8520; // @[digest.scala 81:19 63:25]
  wire  _GEN_9109 = 6'h2a == state ? 1'h0 : _GEN_8603; // @[digest.scala 81:19 68:25]
  wire  _GEN_9192 = 6'h2a == state ? 1'h0 : _GEN_8686; // @[digest.scala 81:19 73:25]
  wire  _GEN_9275 = 6'h2a == state ? 1'h0 : _GEN_8769; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_9276 = 6'h29 == state ? $signed(_t_T_10) : $signed(t); // @[digest.scala 249:15 35:16 81:19]
  wire [5:0] _GEN_9277 = 6'h29 == state ? 6'h2a : _GEN_8771; // @[digest.scala 250:19 81:19]
  wire [31:0] _GEN_9278 = 6'h29 == state ? $signed(e) : $signed(_GEN_8770); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_9279 = 6'h29 == state ? $signed(d) : $signed(_GEN_8772); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_9280 = 6'h29 == state ? $signed(c) : $signed(_GEN_8773); // @[digest.scala 26:16 81:19]
  wire  _GEN_9281 = 6'h29 == state ? 1'h0 : _GEN_8774; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_9284 = 6'h29 == state ? $signed(b) : $signed(_GEN_8777); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_9285 = 6'h29 == state ? $signed(a) : $signed(_GEN_8778); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_9286 = 6'h29 == state ? $signed(j) : $signed(_GEN_8779); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_9287 = 6'h29 == state ? $signed(i) : $signed(_GEN_8780); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_9369 = 6'h29 == state ? $signed(digest_0) : $signed(_GEN_8862); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9370 = 6'h29 == state ? $signed(digest_1) : $signed(_GEN_8863); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9371 = 6'h29 == state ? $signed(digest_2) : $signed(_GEN_8864); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9372 = 6'h29 == state ? $signed(digest_3) : $signed(_GEN_8865); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9373 = 6'h29 == state ? $signed(digest_4) : $signed(_GEN_8866); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9374 = 6'h29 == state ? $signed(digest_5) : $signed(_GEN_8867); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9375 = 6'h29 == state ? $signed(digest_6) : $signed(_GEN_8868); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9376 = 6'h29 == state ? $signed(digest_7) : $signed(_GEN_8869); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9377 = 6'h29 == state ? $signed(digest_8) : $signed(_GEN_8870); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9378 = 6'h29 == state ? $signed(digest_9) : $signed(_GEN_8871); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9379 = 6'h29 == state ? $signed(digest_10) : $signed(_GEN_8872); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9380 = 6'h29 == state ? $signed(digest_11) : $signed(_GEN_8873); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9381 = 6'h29 == state ? $signed(digest_12) : $signed(_GEN_8874); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9382 = 6'h29 == state ? $signed(digest_13) : $signed(_GEN_8875); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9383 = 6'h29 == state ? $signed(digest_14) : $signed(_GEN_8876); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9384 = 6'h29 == state ? $signed(digest_15) : $signed(_GEN_8877); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9385 = 6'h29 == state ? $signed(digest_16) : $signed(_GEN_8878); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9386 = 6'h29 == state ? $signed(digest_17) : $signed(_GEN_8879); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9387 = 6'h29 == state ? $signed(digest_18) : $signed(_GEN_8880); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9388 = 6'h29 == state ? $signed(digest_19) : $signed(_GEN_8881); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9389 = 6'h29 == state ? $signed(digest_20) : $signed(_GEN_8882); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9390 = 6'h29 == state ? $signed(digest_21) : $signed(_GEN_8883); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9391 = 6'h29 == state ? $signed(digest_22) : $signed(_GEN_8884); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9392 = 6'h29 == state ? $signed(digest_23) : $signed(_GEN_8885); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9393 = 6'h29 == state ? $signed(digest_24) : $signed(_GEN_8886); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9394 = 6'h29 == state ? $signed(digest_25) : $signed(_GEN_8887); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9395 = 6'h29 == state ? $signed(digest_26) : $signed(_GEN_8888); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9396 = 6'h29 == state ? $signed(digest_27) : $signed(_GEN_8889); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9397 = 6'h29 == state ? $signed(digest_28) : $signed(_GEN_8890); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9398 = 6'h29 == state ? $signed(digest_29) : $signed(_GEN_8891); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9399 = 6'h29 == state ? $signed(digest_30) : $signed(_GEN_8892); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9400 = 6'h29 == state ? $signed(digest_31) : $signed(_GEN_8893); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9401 = 6'h29 == state ? $signed(digest_32) : $signed(_GEN_8894); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9402 = 6'h29 == state ? $signed(digest_33) : $signed(_GEN_8895); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9403 = 6'h29 == state ? $signed(digest_34) : $signed(_GEN_8896); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9404 = 6'h29 == state ? $signed(digest_35) : $signed(_GEN_8897); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9405 = 6'h29 == state ? $signed(digest_36) : $signed(_GEN_8898); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9406 = 6'h29 == state ? $signed(digest_37) : $signed(_GEN_8899); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9407 = 6'h29 == state ? $signed(digest_38) : $signed(_GEN_8900); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9408 = 6'h29 == state ? $signed(digest_39) : $signed(_GEN_8901); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9409 = 6'h29 == state ? $signed(digest_40) : $signed(_GEN_8902); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9410 = 6'h29 == state ? $signed(digest_41) : $signed(_GEN_8903); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9411 = 6'h29 == state ? $signed(digest_42) : $signed(_GEN_8904); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9412 = 6'h29 == state ? $signed(digest_43) : $signed(_GEN_8905); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9413 = 6'h29 == state ? $signed(digest_44) : $signed(_GEN_8906); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9414 = 6'h29 == state ? $signed(digest_45) : $signed(_GEN_8907); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9415 = 6'h29 == state ? $signed(digest_46) : $signed(_GEN_8908); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9416 = 6'h29 == state ? $signed(digest_47) : $signed(_GEN_8909); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9417 = 6'h29 == state ? $signed(digest_48) : $signed(_GEN_8910); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9418 = 6'h29 == state ? $signed(digest_49) : $signed(_GEN_8911); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9419 = 6'h29 == state ? $signed(digest_50) : $signed(_GEN_8912); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9420 = 6'h29 == state ? $signed(digest_51) : $signed(_GEN_8913); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9421 = 6'h29 == state ? $signed(digest_52) : $signed(_GEN_8914); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9422 = 6'h29 == state ? $signed(digest_53) : $signed(_GEN_8915); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9423 = 6'h29 == state ? $signed(digest_54) : $signed(_GEN_8916); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9424 = 6'h29 == state ? $signed(digest_55) : $signed(_GEN_8917); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9425 = 6'h29 == state ? $signed(digest_56) : $signed(_GEN_8918); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9426 = 6'h29 == state ? $signed(digest_57) : $signed(_GEN_8919); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9427 = 6'h29 == state ? $signed(digest_58) : $signed(_GEN_8920); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9428 = 6'h29 == state ? $signed(digest_59) : $signed(_GEN_8921); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9429 = 6'h29 == state ? $signed(digest_60) : $signed(_GEN_8922); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9430 = 6'h29 == state ? $signed(digest_61) : $signed(_GEN_8923); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9431 = 6'h29 == state ? $signed(digest_62) : $signed(_GEN_8924); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9432 = 6'h29 == state ? $signed(digest_63) : $signed(_GEN_8925); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9433 = 6'h29 == state ? $signed(digest_64) : $signed(_GEN_8926); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9434 = 6'h29 == state ? $signed(digest_65) : $signed(_GEN_8927); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9435 = 6'h29 == state ? $signed(digest_66) : $signed(_GEN_8928); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9436 = 6'h29 == state ? $signed(digest_67) : $signed(_GEN_8929); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9437 = 6'h29 == state ? $signed(digest_68) : $signed(_GEN_8930); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9438 = 6'h29 == state ? $signed(digest_69) : $signed(_GEN_8931); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9439 = 6'h29 == state ? $signed(digest_70) : $signed(_GEN_8932); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9440 = 6'h29 == state ? $signed(digest_71) : $signed(_GEN_8933); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9441 = 6'h29 == state ? $signed(digest_72) : $signed(_GEN_8934); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9442 = 6'h29 == state ? $signed(digest_73) : $signed(_GEN_8935); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9443 = 6'h29 == state ? $signed(digest_74) : $signed(_GEN_8936); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9444 = 6'h29 == state ? $signed(digest_75) : $signed(_GEN_8937); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9445 = 6'h29 == state ? $signed(digest_76) : $signed(_GEN_8938); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9446 = 6'h29 == state ? $signed(digest_77) : $signed(_GEN_8939); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9447 = 6'h29 == state ? $signed(digest_78) : $signed(_GEN_8940); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9448 = 6'h29 == state ? $signed(digest_79) : $signed(_GEN_8941); // @[digest.scala 81:19 53:21]
  wire  _GEN_9450 = 6'h29 == state ? 1'h0 : _GEN_8943; // @[digest.scala 81:19 58:25]
  wire  _GEN_9533 = 6'h29 == state ? 1'h0 : _GEN_9026; // @[digest.scala 81:19 63:25]
  wire  _GEN_9616 = 6'h29 == state ? 1'h0 : _GEN_9109; // @[digest.scala 81:19 68:25]
  wire  _GEN_9699 = 6'h29 == state ? 1'h0 : _GEN_9192; // @[digest.scala 81:19 73:25]
  wire  _GEN_9782 = 6'h29 == state ? 1'h0 : _GEN_9275; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_9783 = 6'h28 == state ? $signed(__m_rol_1_io_out_rol) : $signed(_GEN_9276); // @[digest.scala 242:15 81:19]
  wire  _GEN_9784 = 6'h28 == state & __m_rol_1_io_valid_T; // @[digest.scala 81:19 243:32 48:24]
  wire [5:0] _GEN_9787 = 6'h28 == state ? _state_T_16 : _GEN_9277; // @[digest.scala 246:19 81:19]
  wire [31:0] _GEN_9788 = 6'h28 == state ? $signed(e) : $signed(_GEN_9278); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_9789 = 6'h28 == state ? $signed(d) : $signed(_GEN_9279); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_9790 = 6'h28 == state ? $signed(c) : $signed(_GEN_9280); // @[digest.scala 26:16 81:19]
  wire  _GEN_9791 = 6'h28 == state ? 1'h0 : _GEN_9281; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_9794 = 6'h28 == state ? $signed(b) : $signed(_GEN_9284); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_9795 = 6'h28 == state ? $signed(a) : $signed(_GEN_9285); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_9796 = 6'h28 == state ? $signed(j) : $signed(_GEN_9286); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_9797 = 6'h28 == state ? $signed(i) : $signed(_GEN_9287); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_9879 = 6'h28 == state ? $signed(digest_0) : $signed(_GEN_9369); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9880 = 6'h28 == state ? $signed(digest_1) : $signed(_GEN_9370); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9881 = 6'h28 == state ? $signed(digest_2) : $signed(_GEN_9371); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9882 = 6'h28 == state ? $signed(digest_3) : $signed(_GEN_9372); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9883 = 6'h28 == state ? $signed(digest_4) : $signed(_GEN_9373); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9884 = 6'h28 == state ? $signed(digest_5) : $signed(_GEN_9374); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9885 = 6'h28 == state ? $signed(digest_6) : $signed(_GEN_9375); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9886 = 6'h28 == state ? $signed(digest_7) : $signed(_GEN_9376); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9887 = 6'h28 == state ? $signed(digest_8) : $signed(_GEN_9377); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9888 = 6'h28 == state ? $signed(digest_9) : $signed(_GEN_9378); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9889 = 6'h28 == state ? $signed(digest_10) : $signed(_GEN_9379); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9890 = 6'h28 == state ? $signed(digest_11) : $signed(_GEN_9380); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9891 = 6'h28 == state ? $signed(digest_12) : $signed(_GEN_9381); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9892 = 6'h28 == state ? $signed(digest_13) : $signed(_GEN_9382); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9893 = 6'h28 == state ? $signed(digest_14) : $signed(_GEN_9383); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9894 = 6'h28 == state ? $signed(digest_15) : $signed(_GEN_9384); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9895 = 6'h28 == state ? $signed(digest_16) : $signed(_GEN_9385); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9896 = 6'h28 == state ? $signed(digest_17) : $signed(_GEN_9386); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9897 = 6'h28 == state ? $signed(digest_18) : $signed(_GEN_9387); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9898 = 6'h28 == state ? $signed(digest_19) : $signed(_GEN_9388); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9899 = 6'h28 == state ? $signed(digest_20) : $signed(_GEN_9389); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9900 = 6'h28 == state ? $signed(digest_21) : $signed(_GEN_9390); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9901 = 6'h28 == state ? $signed(digest_22) : $signed(_GEN_9391); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9902 = 6'h28 == state ? $signed(digest_23) : $signed(_GEN_9392); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9903 = 6'h28 == state ? $signed(digest_24) : $signed(_GEN_9393); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9904 = 6'h28 == state ? $signed(digest_25) : $signed(_GEN_9394); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9905 = 6'h28 == state ? $signed(digest_26) : $signed(_GEN_9395); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9906 = 6'h28 == state ? $signed(digest_27) : $signed(_GEN_9396); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9907 = 6'h28 == state ? $signed(digest_28) : $signed(_GEN_9397); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9908 = 6'h28 == state ? $signed(digest_29) : $signed(_GEN_9398); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9909 = 6'h28 == state ? $signed(digest_30) : $signed(_GEN_9399); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9910 = 6'h28 == state ? $signed(digest_31) : $signed(_GEN_9400); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9911 = 6'h28 == state ? $signed(digest_32) : $signed(_GEN_9401); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9912 = 6'h28 == state ? $signed(digest_33) : $signed(_GEN_9402); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9913 = 6'h28 == state ? $signed(digest_34) : $signed(_GEN_9403); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9914 = 6'h28 == state ? $signed(digest_35) : $signed(_GEN_9404); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9915 = 6'h28 == state ? $signed(digest_36) : $signed(_GEN_9405); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9916 = 6'h28 == state ? $signed(digest_37) : $signed(_GEN_9406); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9917 = 6'h28 == state ? $signed(digest_38) : $signed(_GEN_9407); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9918 = 6'h28 == state ? $signed(digest_39) : $signed(_GEN_9408); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9919 = 6'h28 == state ? $signed(digest_40) : $signed(_GEN_9409); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9920 = 6'h28 == state ? $signed(digest_41) : $signed(_GEN_9410); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9921 = 6'h28 == state ? $signed(digest_42) : $signed(_GEN_9411); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9922 = 6'h28 == state ? $signed(digest_43) : $signed(_GEN_9412); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9923 = 6'h28 == state ? $signed(digest_44) : $signed(_GEN_9413); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9924 = 6'h28 == state ? $signed(digest_45) : $signed(_GEN_9414); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9925 = 6'h28 == state ? $signed(digest_46) : $signed(_GEN_9415); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9926 = 6'h28 == state ? $signed(digest_47) : $signed(_GEN_9416); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9927 = 6'h28 == state ? $signed(digest_48) : $signed(_GEN_9417); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9928 = 6'h28 == state ? $signed(digest_49) : $signed(_GEN_9418); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9929 = 6'h28 == state ? $signed(digest_50) : $signed(_GEN_9419); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9930 = 6'h28 == state ? $signed(digest_51) : $signed(_GEN_9420); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9931 = 6'h28 == state ? $signed(digest_52) : $signed(_GEN_9421); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9932 = 6'h28 == state ? $signed(digest_53) : $signed(_GEN_9422); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9933 = 6'h28 == state ? $signed(digest_54) : $signed(_GEN_9423); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9934 = 6'h28 == state ? $signed(digest_55) : $signed(_GEN_9424); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9935 = 6'h28 == state ? $signed(digest_56) : $signed(_GEN_9425); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9936 = 6'h28 == state ? $signed(digest_57) : $signed(_GEN_9426); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9937 = 6'h28 == state ? $signed(digest_58) : $signed(_GEN_9427); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9938 = 6'h28 == state ? $signed(digest_59) : $signed(_GEN_9428); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9939 = 6'h28 == state ? $signed(digest_60) : $signed(_GEN_9429); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9940 = 6'h28 == state ? $signed(digest_61) : $signed(_GEN_9430); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9941 = 6'h28 == state ? $signed(digest_62) : $signed(_GEN_9431); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9942 = 6'h28 == state ? $signed(digest_63) : $signed(_GEN_9432); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9943 = 6'h28 == state ? $signed(digest_64) : $signed(_GEN_9433); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9944 = 6'h28 == state ? $signed(digest_65) : $signed(_GEN_9434); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9945 = 6'h28 == state ? $signed(digest_66) : $signed(_GEN_9435); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9946 = 6'h28 == state ? $signed(digest_67) : $signed(_GEN_9436); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9947 = 6'h28 == state ? $signed(digest_68) : $signed(_GEN_9437); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9948 = 6'h28 == state ? $signed(digest_69) : $signed(_GEN_9438); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9949 = 6'h28 == state ? $signed(digest_70) : $signed(_GEN_9439); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9950 = 6'h28 == state ? $signed(digest_71) : $signed(_GEN_9440); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9951 = 6'h28 == state ? $signed(digest_72) : $signed(_GEN_9441); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9952 = 6'h28 == state ? $signed(digest_73) : $signed(_GEN_9442); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9953 = 6'h28 == state ? $signed(digest_74) : $signed(_GEN_9443); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9954 = 6'h28 == state ? $signed(digest_75) : $signed(_GEN_9444); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9955 = 6'h28 == state ? $signed(digest_76) : $signed(_GEN_9445); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9956 = 6'h28 == state ? $signed(digest_77) : $signed(_GEN_9446); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9957 = 6'h28 == state ? $signed(digest_78) : $signed(_GEN_9447); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_9958 = 6'h28 == state ? $signed(digest_79) : $signed(_GEN_9448); // @[digest.scala 81:19 53:21]
  wire  _GEN_9960 = 6'h28 == state ? 1'h0 : _GEN_9450; // @[digest.scala 81:19 58:25]
  wire  _GEN_10043 = 6'h28 == state ? 1'h0 : _GEN_9533; // @[digest.scala 81:19 63:25]
  wire  _GEN_10126 = 6'h28 == state ? 1'h0 : _GEN_9616; // @[digest.scala 81:19 68:25]
  wire  _GEN_10209 = 6'h28 == state ? 1'h0 : _GEN_9699; // @[digest.scala 81:19 73:25]
  wire  _GEN_10292 = 6'h28 == state ? 1'h0 : _GEN_9782; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_10293 = 6'h27 == state ? $signed(_temp_T_81) : $signed(temp); // @[digest.scala 238:18 38:19 81:19]
  wire [5:0] _GEN_10294 = 6'h27 == state ? 6'h28 : _GEN_9787; // @[digest.scala 239:19 81:19]
  wire [31:0] _GEN_10295 = 6'h27 == state ? $signed(t) : $signed(_GEN_9783); // @[digest.scala 35:16 81:19]
  wire  _GEN_10296 = 6'h27 == state ? 1'h0 : _GEN_9784; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_10299 = 6'h27 == state ? $signed(e) : $signed(_GEN_9788); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_10300 = 6'h27 == state ? $signed(d) : $signed(_GEN_9789); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_10301 = 6'h27 == state ? $signed(c) : $signed(_GEN_9790); // @[digest.scala 26:16 81:19]
  wire  _GEN_10302 = 6'h27 == state ? 1'h0 : _GEN_9791; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_10305 = 6'h27 == state ? $signed(b) : $signed(_GEN_9794); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_10306 = 6'h27 == state ? $signed(a) : $signed(_GEN_9795); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_10307 = 6'h27 == state ? $signed(j) : $signed(_GEN_9796); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_10308 = 6'h27 == state ? $signed(i) : $signed(_GEN_9797); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_10390 = 6'h27 == state ? $signed(digest_0) : $signed(_GEN_9879); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10391 = 6'h27 == state ? $signed(digest_1) : $signed(_GEN_9880); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10392 = 6'h27 == state ? $signed(digest_2) : $signed(_GEN_9881); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10393 = 6'h27 == state ? $signed(digest_3) : $signed(_GEN_9882); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10394 = 6'h27 == state ? $signed(digest_4) : $signed(_GEN_9883); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10395 = 6'h27 == state ? $signed(digest_5) : $signed(_GEN_9884); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10396 = 6'h27 == state ? $signed(digest_6) : $signed(_GEN_9885); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10397 = 6'h27 == state ? $signed(digest_7) : $signed(_GEN_9886); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10398 = 6'h27 == state ? $signed(digest_8) : $signed(_GEN_9887); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10399 = 6'h27 == state ? $signed(digest_9) : $signed(_GEN_9888); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10400 = 6'h27 == state ? $signed(digest_10) : $signed(_GEN_9889); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10401 = 6'h27 == state ? $signed(digest_11) : $signed(_GEN_9890); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10402 = 6'h27 == state ? $signed(digest_12) : $signed(_GEN_9891); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10403 = 6'h27 == state ? $signed(digest_13) : $signed(_GEN_9892); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10404 = 6'h27 == state ? $signed(digest_14) : $signed(_GEN_9893); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10405 = 6'h27 == state ? $signed(digest_15) : $signed(_GEN_9894); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10406 = 6'h27 == state ? $signed(digest_16) : $signed(_GEN_9895); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10407 = 6'h27 == state ? $signed(digest_17) : $signed(_GEN_9896); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10408 = 6'h27 == state ? $signed(digest_18) : $signed(_GEN_9897); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10409 = 6'h27 == state ? $signed(digest_19) : $signed(_GEN_9898); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10410 = 6'h27 == state ? $signed(digest_20) : $signed(_GEN_9899); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10411 = 6'h27 == state ? $signed(digest_21) : $signed(_GEN_9900); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10412 = 6'h27 == state ? $signed(digest_22) : $signed(_GEN_9901); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10413 = 6'h27 == state ? $signed(digest_23) : $signed(_GEN_9902); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10414 = 6'h27 == state ? $signed(digest_24) : $signed(_GEN_9903); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10415 = 6'h27 == state ? $signed(digest_25) : $signed(_GEN_9904); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10416 = 6'h27 == state ? $signed(digest_26) : $signed(_GEN_9905); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10417 = 6'h27 == state ? $signed(digest_27) : $signed(_GEN_9906); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10418 = 6'h27 == state ? $signed(digest_28) : $signed(_GEN_9907); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10419 = 6'h27 == state ? $signed(digest_29) : $signed(_GEN_9908); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10420 = 6'h27 == state ? $signed(digest_30) : $signed(_GEN_9909); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10421 = 6'h27 == state ? $signed(digest_31) : $signed(_GEN_9910); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10422 = 6'h27 == state ? $signed(digest_32) : $signed(_GEN_9911); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10423 = 6'h27 == state ? $signed(digest_33) : $signed(_GEN_9912); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10424 = 6'h27 == state ? $signed(digest_34) : $signed(_GEN_9913); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10425 = 6'h27 == state ? $signed(digest_35) : $signed(_GEN_9914); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10426 = 6'h27 == state ? $signed(digest_36) : $signed(_GEN_9915); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10427 = 6'h27 == state ? $signed(digest_37) : $signed(_GEN_9916); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10428 = 6'h27 == state ? $signed(digest_38) : $signed(_GEN_9917); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10429 = 6'h27 == state ? $signed(digest_39) : $signed(_GEN_9918); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10430 = 6'h27 == state ? $signed(digest_40) : $signed(_GEN_9919); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10431 = 6'h27 == state ? $signed(digest_41) : $signed(_GEN_9920); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10432 = 6'h27 == state ? $signed(digest_42) : $signed(_GEN_9921); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10433 = 6'h27 == state ? $signed(digest_43) : $signed(_GEN_9922); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10434 = 6'h27 == state ? $signed(digest_44) : $signed(_GEN_9923); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10435 = 6'h27 == state ? $signed(digest_45) : $signed(_GEN_9924); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10436 = 6'h27 == state ? $signed(digest_46) : $signed(_GEN_9925); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10437 = 6'h27 == state ? $signed(digest_47) : $signed(_GEN_9926); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10438 = 6'h27 == state ? $signed(digest_48) : $signed(_GEN_9927); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10439 = 6'h27 == state ? $signed(digest_49) : $signed(_GEN_9928); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10440 = 6'h27 == state ? $signed(digest_50) : $signed(_GEN_9929); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10441 = 6'h27 == state ? $signed(digest_51) : $signed(_GEN_9930); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10442 = 6'h27 == state ? $signed(digest_52) : $signed(_GEN_9931); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10443 = 6'h27 == state ? $signed(digest_53) : $signed(_GEN_9932); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10444 = 6'h27 == state ? $signed(digest_54) : $signed(_GEN_9933); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10445 = 6'h27 == state ? $signed(digest_55) : $signed(_GEN_9934); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10446 = 6'h27 == state ? $signed(digest_56) : $signed(_GEN_9935); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10447 = 6'h27 == state ? $signed(digest_57) : $signed(_GEN_9936); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10448 = 6'h27 == state ? $signed(digest_58) : $signed(_GEN_9937); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10449 = 6'h27 == state ? $signed(digest_59) : $signed(_GEN_9938); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10450 = 6'h27 == state ? $signed(digest_60) : $signed(_GEN_9939); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10451 = 6'h27 == state ? $signed(digest_61) : $signed(_GEN_9940); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10452 = 6'h27 == state ? $signed(digest_62) : $signed(_GEN_9941); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10453 = 6'h27 == state ? $signed(digest_63) : $signed(_GEN_9942); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10454 = 6'h27 == state ? $signed(digest_64) : $signed(_GEN_9943); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10455 = 6'h27 == state ? $signed(digest_65) : $signed(_GEN_9944); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10456 = 6'h27 == state ? $signed(digest_66) : $signed(_GEN_9945); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10457 = 6'h27 == state ? $signed(digest_67) : $signed(_GEN_9946); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10458 = 6'h27 == state ? $signed(digest_68) : $signed(_GEN_9947); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10459 = 6'h27 == state ? $signed(digest_69) : $signed(_GEN_9948); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10460 = 6'h27 == state ? $signed(digest_70) : $signed(_GEN_9949); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10461 = 6'h27 == state ? $signed(digest_71) : $signed(_GEN_9950); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10462 = 6'h27 == state ? $signed(digest_72) : $signed(_GEN_9951); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10463 = 6'h27 == state ? $signed(digest_73) : $signed(_GEN_9952); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10464 = 6'h27 == state ? $signed(digest_74) : $signed(_GEN_9953); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10465 = 6'h27 == state ? $signed(digest_75) : $signed(_GEN_9954); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10466 = 6'h27 == state ? $signed(digest_76) : $signed(_GEN_9955); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10467 = 6'h27 == state ? $signed(digest_77) : $signed(_GEN_9956); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10468 = 6'h27 == state ? $signed(digest_78) : $signed(_GEN_9957); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10469 = 6'h27 == state ? $signed(digest_79) : $signed(_GEN_9958); // @[digest.scala 81:19 53:21]
  wire  _GEN_10471 = 6'h27 == state ? 1'h0 : _GEN_9960; // @[digest.scala 81:19 58:25]
  wire  _GEN_10554 = 6'h27 == state ? 1'h0 : _GEN_10043; // @[digest.scala 81:19 63:25]
  wire  _GEN_10637 = 6'h27 == state ? 1'h0 : _GEN_10126; // @[digest.scala 81:19 68:25]
  wire  _GEN_10720 = 6'h27 == state ? 1'h0 : _GEN_10209; // @[digest.scala 81:19 73:25]
  wire  _GEN_10803 = 6'h27 == state ? 1'h0 : _GEN_10292; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_10804 = 6'h26 == state ? $signed(_temp_T_58) : $signed(_GEN_10293); // @[digest.scala 234:18 81:19]
  wire [5:0] _GEN_10805 = 6'h26 == state ? 6'h27 : _GEN_10294; // @[digest.scala 235:19 81:19]
  wire [31:0] _GEN_10806 = 6'h26 == state ? $signed(t) : $signed(_GEN_10295); // @[digest.scala 35:16 81:19]
  wire  _GEN_10807 = 6'h26 == state ? 1'h0 : _GEN_10296; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_10810 = 6'h26 == state ? $signed(e) : $signed(_GEN_10299); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_10811 = 6'h26 == state ? $signed(d) : $signed(_GEN_10300); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_10812 = 6'h26 == state ? $signed(c) : $signed(_GEN_10301); // @[digest.scala 26:16 81:19]
  wire  _GEN_10813 = 6'h26 == state ? 1'h0 : _GEN_10302; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_10816 = 6'h26 == state ? $signed(b) : $signed(_GEN_10305); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_10817 = 6'h26 == state ? $signed(a) : $signed(_GEN_10306); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_10818 = 6'h26 == state ? $signed(j) : $signed(_GEN_10307); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_10819 = 6'h26 == state ? $signed(i) : $signed(_GEN_10308); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_10901 = 6'h26 == state ? $signed(digest_0) : $signed(_GEN_10390); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10902 = 6'h26 == state ? $signed(digest_1) : $signed(_GEN_10391); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10903 = 6'h26 == state ? $signed(digest_2) : $signed(_GEN_10392); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10904 = 6'h26 == state ? $signed(digest_3) : $signed(_GEN_10393); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10905 = 6'h26 == state ? $signed(digest_4) : $signed(_GEN_10394); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10906 = 6'h26 == state ? $signed(digest_5) : $signed(_GEN_10395); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10907 = 6'h26 == state ? $signed(digest_6) : $signed(_GEN_10396); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10908 = 6'h26 == state ? $signed(digest_7) : $signed(_GEN_10397); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10909 = 6'h26 == state ? $signed(digest_8) : $signed(_GEN_10398); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10910 = 6'h26 == state ? $signed(digest_9) : $signed(_GEN_10399); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10911 = 6'h26 == state ? $signed(digest_10) : $signed(_GEN_10400); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10912 = 6'h26 == state ? $signed(digest_11) : $signed(_GEN_10401); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10913 = 6'h26 == state ? $signed(digest_12) : $signed(_GEN_10402); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10914 = 6'h26 == state ? $signed(digest_13) : $signed(_GEN_10403); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10915 = 6'h26 == state ? $signed(digest_14) : $signed(_GEN_10404); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10916 = 6'h26 == state ? $signed(digest_15) : $signed(_GEN_10405); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10917 = 6'h26 == state ? $signed(digest_16) : $signed(_GEN_10406); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10918 = 6'h26 == state ? $signed(digest_17) : $signed(_GEN_10407); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10919 = 6'h26 == state ? $signed(digest_18) : $signed(_GEN_10408); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10920 = 6'h26 == state ? $signed(digest_19) : $signed(_GEN_10409); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10921 = 6'h26 == state ? $signed(digest_20) : $signed(_GEN_10410); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10922 = 6'h26 == state ? $signed(digest_21) : $signed(_GEN_10411); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10923 = 6'h26 == state ? $signed(digest_22) : $signed(_GEN_10412); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10924 = 6'h26 == state ? $signed(digest_23) : $signed(_GEN_10413); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10925 = 6'h26 == state ? $signed(digest_24) : $signed(_GEN_10414); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10926 = 6'h26 == state ? $signed(digest_25) : $signed(_GEN_10415); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10927 = 6'h26 == state ? $signed(digest_26) : $signed(_GEN_10416); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10928 = 6'h26 == state ? $signed(digest_27) : $signed(_GEN_10417); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10929 = 6'h26 == state ? $signed(digest_28) : $signed(_GEN_10418); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10930 = 6'h26 == state ? $signed(digest_29) : $signed(_GEN_10419); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10931 = 6'h26 == state ? $signed(digest_30) : $signed(_GEN_10420); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10932 = 6'h26 == state ? $signed(digest_31) : $signed(_GEN_10421); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10933 = 6'h26 == state ? $signed(digest_32) : $signed(_GEN_10422); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10934 = 6'h26 == state ? $signed(digest_33) : $signed(_GEN_10423); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10935 = 6'h26 == state ? $signed(digest_34) : $signed(_GEN_10424); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10936 = 6'h26 == state ? $signed(digest_35) : $signed(_GEN_10425); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10937 = 6'h26 == state ? $signed(digest_36) : $signed(_GEN_10426); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10938 = 6'h26 == state ? $signed(digest_37) : $signed(_GEN_10427); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10939 = 6'h26 == state ? $signed(digest_38) : $signed(_GEN_10428); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10940 = 6'h26 == state ? $signed(digest_39) : $signed(_GEN_10429); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10941 = 6'h26 == state ? $signed(digest_40) : $signed(_GEN_10430); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10942 = 6'h26 == state ? $signed(digest_41) : $signed(_GEN_10431); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10943 = 6'h26 == state ? $signed(digest_42) : $signed(_GEN_10432); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10944 = 6'h26 == state ? $signed(digest_43) : $signed(_GEN_10433); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10945 = 6'h26 == state ? $signed(digest_44) : $signed(_GEN_10434); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10946 = 6'h26 == state ? $signed(digest_45) : $signed(_GEN_10435); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10947 = 6'h26 == state ? $signed(digest_46) : $signed(_GEN_10436); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10948 = 6'h26 == state ? $signed(digest_47) : $signed(_GEN_10437); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10949 = 6'h26 == state ? $signed(digest_48) : $signed(_GEN_10438); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10950 = 6'h26 == state ? $signed(digest_49) : $signed(_GEN_10439); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10951 = 6'h26 == state ? $signed(digest_50) : $signed(_GEN_10440); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10952 = 6'h26 == state ? $signed(digest_51) : $signed(_GEN_10441); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10953 = 6'h26 == state ? $signed(digest_52) : $signed(_GEN_10442); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10954 = 6'h26 == state ? $signed(digest_53) : $signed(_GEN_10443); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10955 = 6'h26 == state ? $signed(digest_54) : $signed(_GEN_10444); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10956 = 6'h26 == state ? $signed(digest_55) : $signed(_GEN_10445); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10957 = 6'h26 == state ? $signed(digest_56) : $signed(_GEN_10446); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10958 = 6'h26 == state ? $signed(digest_57) : $signed(_GEN_10447); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10959 = 6'h26 == state ? $signed(digest_58) : $signed(_GEN_10448); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10960 = 6'h26 == state ? $signed(digest_59) : $signed(_GEN_10449); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10961 = 6'h26 == state ? $signed(digest_60) : $signed(_GEN_10450); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10962 = 6'h26 == state ? $signed(digest_61) : $signed(_GEN_10451); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10963 = 6'h26 == state ? $signed(digest_62) : $signed(_GEN_10452); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10964 = 6'h26 == state ? $signed(digest_63) : $signed(_GEN_10453); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10965 = 6'h26 == state ? $signed(digest_64) : $signed(_GEN_10454); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10966 = 6'h26 == state ? $signed(digest_65) : $signed(_GEN_10455); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10967 = 6'h26 == state ? $signed(digest_66) : $signed(_GEN_10456); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10968 = 6'h26 == state ? $signed(digest_67) : $signed(_GEN_10457); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10969 = 6'h26 == state ? $signed(digest_68) : $signed(_GEN_10458); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10970 = 6'h26 == state ? $signed(digest_69) : $signed(_GEN_10459); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10971 = 6'h26 == state ? $signed(digest_70) : $signed(_GEN_10460); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10972 = 6'h26 == state ? $signed(digest_71) : $signed(_GEN_10461); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10973 = 6'h26 == state ? $signed(digest_72) : $signed(_GEN_10462); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10974 = 6'h26 == state ? $signed(digest_73) : $signed(_GEN_10463); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10975 = 6'h26 == state ? $signed(digest_74) : $signed(_GEN_10464); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10976 = 6'h26 == state ? $signed(digest_75) : $signed(_GEN_10465); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10977 = 6'h26 == state ? $signed(digest_76) : $signed(_GEN_10466); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10978 = 6'h26 == state ? $signed(digest_77) : $signed(_GEN_10467); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10979 = 6'h26 == state ? $signed(digest_78) : $signed(_GEN_10468); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_10980 = 6'h26 == state ? $signed(digest_79) : $signed(_GEN_10469); // @[digest.scala 81:19 53:21]
  wire  _GEN_10982 = 6'h26 == state ? 1'h0 : _GEN_10471; // @[digest.scala 81:19 58:25]
  wire  _GEN_11065 = 6'h26 == state ? 1'h0 : _GEN_10554; // @[digest.scala 81:19 63:25]
  wire  _GEN_11148 = 6'h26 == state ? 1'h0 : _GEN_10637; // @[digest.scala 81:19 68:25]
  wire  _GEN_11231 = 6'h26 == state ? 1'h0 : _GEN_10720; // @[digest.scala 81:19 73:25]
  wire  _GEN_11314 = 6'h26 == state ? 1'h0 : _GEN_10803; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_11315 = 6'h25 == state ? $signed(_temp_T_74) : $signed(_GEN_10804); // @[digest.scala 230:18 81:19]
  wire [5:0] _GEN_11316 = 6'h25 == state ? 6'h28 : _GEN_10805; // @[digest.scala 231:19 81:19]
  wire [31:0] _GEN_11317 = 6'h25 == state ? $signed(t) : $signed(_GEN_10806); // @[digest.scala 35:16 81:19]
  wire  _GEN_11318 = 6'h25 == state ? 1'h0 : _GEN_10807; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_11321 = 6'h25 == state ? $signed(e) : $signed(_GEN_10810); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_11322 = 6'h25 == state ? $signed(d) : $signed(_GEN_10811); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_11323 = 6'h25 == state ? $signed(c) : $signed(_GEN_10812); // @[digest.scala 26:16 81:19]
  wire  _GEN_11324 = 6'h25 == state ? 1'h0 : _GEN_10813; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_11327 = 6'h25 == state ? $signed(b) : $signed(_GEN_10816); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_11328 = 6'h25 == state ? $signed(a) : $signed(_GEN_10817); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_11329 = 6'h25 == state ? $signed(j) : $signed(_GEN_10818); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_11330 = 6'h25 == state ? $signed(i) : $signed(_GEN_10819); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_11412 = 6'h25 == state ? $signed(digest_0) : $signed(_GEN_10901); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11413 = 6'h25 == state ? $signed(digest_1) : $signed(_GEN_10902); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11414 = 6'h25 == state ? $signed(digest_2) : $signed(_GEN_10903); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11415 = 6'h25 == state ? $signed(digest_3) : $signed(_GEN_10904); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11416 = 6'h25 == state ? $signed(digest_4) : $signed(_GEN_10905); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11417 = 6'h25 == state ? $signed(digest_5) : $signed(_GEN_10906); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11418 = 6'h25 == state ? $signed(digest_6) : $signed(_GEN_10907); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11419 = 6'h25 == state ? $signed(digest_7) : $signed(_GEN_10908); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11420 = 6'h25 == state ? $signed(digest_8) : $signed(_GEN_10909); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11421 = 6'h25 == state ? $signed(digest_9) : $signed(_GEN_10910); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11422 = 6'h25 == state ? $signed(digest_10) : $signed(_GEN_10911); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11423 = 6'h25 == state ? $signed(digest_11) : $signed(_GEN_10912); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11424 = 6'h25 == state ? $signed(digest_12) : $signed(_GEN_10913); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11425 = 6'h25 == state ? $signed(digest_13) : $signed(_GEN_10914); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11426 = 6'h25 == state ? $signed(digest_14) : $signed(_GEN_10915); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11427 = 6'h25 == state ? $signed(digest_15) : $signed(_GEN_10916); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11428 = 6'h25 == state ? $signed(digest_16) : $signed(_GEN_10917); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11429 = 6'h25 == state ? $signed(digest_17) : $signed(_GEN_10918); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11430 = 6'h25 == state ? $signed(digest_18) : $signed(_GEN_10919); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11431 = 6'h25 == state ? $signed(digest_19) : $signed(_GEN_10920); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11432 = 6'h25 == state ? $signed(digest_20) : $signed(_GEN_10921); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11433 = 6'h25 == state ? $signed(digest_21) : $signed(_GEN_10922); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11434 = 6'h25 == state ? $signed(digest_22) : $signed(_GEN_10923); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11435 = 6'h25 == state ? $signed(digest_23) : $signed(_GEN_10924); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11436 = 6'h25 == state ? $signed(digest_24) : $signed(_GEN_10925); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11437 = 6'h25 == state ? $signed(digest_25) : $signed(_GEN_10926); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11438 = 6'h25 == state ? $signed(digest_26) : $signed(_GEN_10927); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11439 = 6'h25 == state ? $signed(digest_27) : $signed(_GEN_10928); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11440 = 6'h25 == state ? $signed(digest_28) : $signed(_GEN_10929); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11441 = 6'h25 == state ? $signed(digest_29) : $signed(_GEN_10930); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11442 = 6'h25 == state ? $signed(digest_30) : $signed(_GEN_10931); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11443 = 6'h25 == state ? $signed(digest_31) : $signed(_GEN_10932); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11444 = 6'h25 == state ? $signed(digest_32) : $signed(_GEN_10933); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11445 = 6'h25 == state ? $signed(digest_33) : $signed(_GEN_10934); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11446 = 6'h25 == state ? $signed(digest_34) : $signed(_GEN_10935); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11447 = 6'h25 == state ? $signed(digest_35) : $signed(_GEN_10936); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11448 = 6'h25 == state ? $signed(digest_36) : $signed(_GEN_10937); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11449 = 6'h25 == state ? $signed(digest_37) : $signed(_GEN_10938); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11450 = 6'h25 == state ? $signed(digest_38) : $signed(_GEN_10939); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11451 = 6'h25 == state ? $signed(digest_39) : $signed(_GEN_10940); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11452 = 6'h25 == state ? $signed(digest_40) : $signed(_GEN_10941); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11453 = 6'h25 == state ? $signed(digest_41) : $signed(_GEN_10942); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11454 = 6'h25 == state ? $signed(digest_42) : $signed(_GEN_10943); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11455 = 6'h25 == state ? $signed(digest_43) : $signed(_GEN_10944); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11456 = 6'h25 == state ? $signed(digest_44) : $signed(_GEN_10945); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11457 = 6'h25 == state ? $signed(digest_45) : $signed(_GEN_10946); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11458 = 6'h25 == state ? $signed(digest_46) : $signed(_GEN_10947); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11459 = 6'h25 == state ? $signed(digest_47) : $signed(_GEN_10948); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11460 = 6'h25 == state ? $signed(digest_48) : $signed(_GEN_10949); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11461 = 6'h25 == state ? $signed(digest_49) : $signed(_GEN_10950); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11462 = 6'h25 == state ? $signed(digest_50) : $signed(_GEN_10951); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11463 = 6'h25 == state ? $signed(digest_51) : $signed(_GEN_10952); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11464 = 6'h25 == state ? $signed(digest_52) : $signed(_GEN_10953); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11465 = 6'h25 == state ? $signed(digest_53) : $signed(_GEN_10954); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11466 = 6'h25 == state ? $signed(digest_54) : $signed(_GEN_10955); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11467 = 6'h25 == state ? $signed(digest_55) : $signed(_GEN_10956); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11468 = 6'h25 == state ? $signed(digest_56) : $signed(_GEN_10957); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11469 = 6'h25 == state ? $signed(digest_57) : $signed(_GEN_10958); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11470 = 6'h25 == state ? $signed(digest_58) : $signed(_GEN_10959); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11471 = 6'h25 == state ? $signed(digest_59) : $signed(_GEN_10960); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11472 = 6'h25 == state ? $signed(digest_60) : $signed(_GEN_10961); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11473 = 6'h25 == state ? $signed(digest_61) : $signed(_GEN_10962); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11474 = 6'h25 == state ? $signed(digest_62) : $signed(_GEN_10963); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11475 = 6'h25 == state ? $signed(digest_63) : $signed(_GEN_10964); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11476 = 6'h25 == state ? $signed(digest_64) : $signed(_GEN_10965); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11477 = 6'h25 == state ? $signed(digest_65) : $signed(_GEN_10966); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11478 = 6'h25 == state ? $signed(digest_66) : $signed(_GEN_10967); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11479 = 6'h25 == state ? $signed(digest_67) : $signed(_GEN_10968); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11480 = 6'h25 == state ? $signed(digest_68) : $signed(_GEN_10969); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11481 = 6'h25 == state ? $signed(digest_69) : $signed(_GEN_10970); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11482 = 6'h25 == state ? $signed(digest_70) : $signed(_GEN_10971); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11483 = 6'h25 == state ? $signed(digest_71) : $signed(_GEN_10972); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11484 = 6'h25 == state ? $signed(digest_72) : $signed(_GEN_10973); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11485 = 6'h25 == state ? $signed(digest_73) : $signed(_GEN_10974); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11486 = 6'h25 == state ? $signed(digest_74) : $signed(_GEN_10975); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11487 = 6'h25 == state ? $signed(digest_75) : $signed(_GEN_10976); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11488 = 6'h25 == state ? $signed(digest_76) : $signed(_GEN_10977); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11489 = 6'h25 == state ? $signed(digest_77) : $signed(_GEN_10978); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11490 = 6'h25 == state ? $signed(digest_78) : $signed(_GEN_10979); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11491 = 6'h25 == state ? $signed(digest_79) : $signed(_GEN_10980); // @[digest.scala 81:19 53:21]
  wire  _GEN_11493 = 6'h25 == state ? 1'h0 : _GEN_10982; // @[digest.scala 81:19 58:25]
  wire  _GEN_11576 = 6'h25 == state ? 1'h0 : _GEN_11065; // @[digest.scala 81:19 63:25]
  wire  _GEN_11659 = 6'h25 == state ? 1'h0 : _GEN_11148; // @[digest.scala 81:19 68:25]
  wire  _GEN_11742 = 6'h25 == state ? 1'h0 : _GEN_11231; // @[digest.scala 81:19 73:25]
  wire  _GEN_11825 = 6'h25 == state ? 1'h0 : _GEN_11314; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_11826 = 6'h24 == state ? $signed(_temp_T_71) : $signed(_GEN_11315); // @[digest.scala 226:18 81:19]
  wire [5:0] _GEN_11827 = 6'h24 == state ? 6'h25 : _GEN_11316; // @[digest.scala 227:19 81:19]
  wire [31:0] _GEN_11828 = 6'h24 == state ? $signed(t) : $signed(_GEN_11317); // @[digest.scala 35:16 81:19]
  wire  _GEN_11829 = 6'h24 == state ? 1'h0 : _GEN_11318; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_11832 = 6'h24 == state ? $signed(e) : $signed(_GEN_11321); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_11833 = 6'h24 == state ? $signed(d) : $signed(_GEN_11322); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_11834 = 6'h24 == state ? $signed(c) : $signed(_GEN_11323); // @[digest.scala 26:16 81:19]
  wire  _GEN_11835 = 6'h24 == state ? 1'h0 : _GEN_11324; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_11838 = 6'h24 == state ? $signed(b) : $signed(_GEN_11327); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_11839 = 6'h24 == state ? $signed(a) : $signed(_GEN_11328); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_11840 = 6'h24 == state ? $signed(j) : $signed(_GEN_11329); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_11841 = 6'h24 == state ? $signed(i) : $signed(_GEN_11330); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_11923 = 6'h24 == state ? $signed(digest_0) : $signed(_GEN_11412); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11924 = 6'h24 == state ? $signed(digest_1) : $signed(_GEN_11413); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11925 = 6'h24 == state ? $signed(digest_2) : $signed(_GEN_11414); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11926 = 6'h24 == state ? $signed(digest_3) : $signed(_GEN_11415); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11927 = 6'h24 == state ? $signed(digest_4) : $signed(_GEN_11416); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11928 = 6'h24 == state ? $signed(digest_5) : $signed(_GEN_11417); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11929 = 6'h24 == state ? $signed(digest_6) : $signed(_GEN_11418); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11930 = 6'h24 == state ? $signed(digest_7) : $signed(_GEN_11419); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11931 = 6'h24 == state ? $signed(digest_8) : $signed(_GEN_11420); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11932 = 6'h24 == state ? $signed(digest_9) : $signed(_GEN_11421); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11933 = 6'h24 == state ? $signed(digest_10) : $signed(_GEN_11422); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11934 = 6'h24 == state ? $signed(digest_11) : $signed(_GEN_11423); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11935 = 6'h24 == state ? $signed(digest_12) : $signed(_GEN_11424); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11936 = 6'h24 == state ? $signed(digest_13) : $signed(_GEN_11425); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11937 = 6'h24 == state ? $signed(digest_14) : $signed(_GEN_11426); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11938 = 6'h24 == state ? $signed(digest_15) : $signed(_GEN_11427); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11939 = 6'h24 == state ? $signed(digest_16) : $signed(_GEN_11428); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11940 = 6'h24 == state ? $signed(digest_17) : $signed(_GEN_11429); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11941 = 6'h24 == state ? $signed(digest_18) : $signed(_GEN_11430); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11942 = 6'h24 == state ? $signed(digest_19) : $signed(_GEN_11431); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11943 = 6'h24 == state ? $signed(digest_20) : $signed(_GEN_11432); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11944 = 6'h24 == state ? $signed(digest_21) : $signed(_GEN_11433); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11945 = 6'h24 == state ? $signed(digest_22) : $signed(_GEN_11434); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11946 = 6'h24 == state ? $signed(digest_23) : $signed(_GEN_11435); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11947 = 6'h24 == state ? $signed(digest_24) : $signed(_GEN_11436); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11948 = 6'h24 == state ? $signed(digest_25) : $signed(_GEN_11437); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11949 = 6'h24 == state ? $signed(digest_26) : $signed(_GEN_11438); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11950 = 6'h24 == state ? $signed(digest_27) : $signed(_GEN_11439); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11951 = 6'h24 == state ? $signed(digest_28) : $signed(_GEN_11440); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11952 = 6'h24 == state ? $signed(digest_29) : $signed(_GEN_11441); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11953 = 6'h24 == state ? $signed(digest_30) : $signed(_GEN_11442); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11954 = 6'h24 == state ? $signed(digest_31) : $signed(_GEN_11443); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11955 = 6'h24 == state ? $signed(digest_32) : $signed(_GEN_11444); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11956 = 6'h24 == state ? $signed(digest_33) : $signed(_GEN_11445); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11957 = 6'h24 == state ? $signed(digest_34) : $signed(_GEN_11446); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11958 = 6'h24 == state ? $signed(digest_35) : $signed(_GEN_11447); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11959 = 6'h24 == state ? $signed(digest_36) : $signed(_GEN_11448); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11960 = 6'h24 == state ? $signed(digest_37) : $signed(_GEN_11449); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11961 = 6'h24 == state ? $signed(digest_38) : $signed(_GEN_11450); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11962 = 6'h24 == state ? $signed(digest_39) : $signed(_GEN_11451); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11963 = 6'h24 == state ? $signed(digest_40) : $signed(_GEN_11452); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11964 = 6'h24 == state ? $signed(digest_41) : $signed(_GEN_11453); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11965 = 6'h24 == state ? $signed(digest_42) : $signed(_GEN_11454); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11966 = 6'h24 == state ? $signed(digest_43) : $signed(_GEN_11455); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11967 = 6'h24 == state ? $signed(digest_44) : $signed(_GEN_11456); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11968 = 6'h24 == state ? $signed(digest_45) : $signed(_GEN_11457); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11969 = 6'h24 == state ? $signed(digest_46) : $signed(_GEN_11458); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11970 = 6'h24 == state ? $signed(digest_47) : $signed(_GEN_11459); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11971 = 6'h24 == state ? $signed(digest_48) : $signed(_GEN_11460); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11972 = 6'h24 == state ? $signed(digest_49) : $signed(_GEN_11461); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11973 = 6'h24 == state ? $signed(digest_50) : $signed(_GEN_11462); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11974 = 6'h24 == state ? $signed(digest_51) : $signed(_GEN_11463); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11975 = 6'h24 == state ? $signed(digest_52) : $signed(_GEN_11464); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11976 = 6'h24 == state ? $signed(digest_53) : $signed(_GEN_11465); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11977 = 6'h24 == state ? $signed(digest_54) : $signed(_GEN_11466); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11978 = 6'h24 == state ? $signed(digest_55) : $signed(_GEN_11467); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11979 = 6'h24 == state ? $signed(digest_56) : $signed(_GEN_11468); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11980 = 6'h24 == state ? $signed(digest_57) : $signed(_GEN_11469); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11981 = 6'h24 == state ? $signed(digest_58) : $signed(_GEN_11470); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11982 = 6'h24 == state ? $signed(digest_59) : $signed(_GEN_11471); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11983 = 6'h24 == state ? $signed(digest_60) : $signed(_GEN_11472); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11984 = 6'h24 == state ? $signed(digest_61) : $signed(_GEN_11473); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11985 = 6'h24 == state ? $signed(digest_62) : $signed(_GEN_11474); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11986 = 6'h24 == state ? $signed(digest_63) : $signed(_GEN_11475); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11987 = 6'h24 == state ? $signed(digest_64) : $signed(_GEN_11476); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11988 = 6'h24 == state ? $signed(digest_65) : $signed(_GEN_11477); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11989 = 6'h24 == state ? $signed(digest_66) : $signed(_GEN_11478); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11990 = 6'h24 == state ? $signed(digest_67) : $signed(_GEN_11479); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11991 = 6'h24 == state ? $signed(digest_68) : $signed(_GEN_11480); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11992 = 6'h24 == state ? $signed(digest_69) : $signed(_GEN_11481); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11993 = 6'h24 == state ? $signed(digest_70) : $signed(_GEN_11482); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11994 = 6'h24 == state ? $signed(digest_71) : $signed(_GEN_11483); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11995 = 6'h24 == state ? $signed(digest_72) : $signed(_GEN_11484); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11996 = 6'h24 == state ? $signed(digest_73) : $signed(_GEN_11485); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11997 = 6'h24 == state ? $signed(digest_74) : $signed(_GEN_11486); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11998 = 6'h24 == state ? $signed(digest_75) : $signed(_GEN_11487); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_11999 = 6'h24 == state ? $signed(digest_76) : $signed(_GEN_11488); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12000 = 6'h24 == state ? $signed(digest_77) : $signed(_GEN_11489); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12001 = 6'h24 == state ? $signed(digest_78) : $signed(_GEN_11490); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12002 = 6'h24 == state ? $signed(digest_79) : $signed(_GEN_11491); // @[digest.scala 81:19 53:21]
  wire  _GEN_12004 = 6'h24 == state ? 1'h0 : _GEN_11493; // @[digest.scala 81:19 58:25]
  wire  _GEN_12087 = 6'h24 == state ? 1'h0 : _GEN_11576; // @[digest.scala 81:19 63:25]
  wire  _GEN_12170 = 6'h24 == state ? 1'h0 : _GEN_11659; // @[digest.scala 81:19 68:25]
  wire  _GEN_12253 = 6'h24 == state ? 1'h0 : _GEN_11742; // @[digest.scala 81:19 73:25]
  wire  _GEN_12336 = 6'h24 == state ? 1'h0 : _GEN_11825; // @[digest.scala 81:19 78:25]
  wire [5:0] _GEN_12337 = 6'h23 == state ? _state_T_15 : _GEN_11827; // @[digest.scala 223:19 81:19]
  wire [31:0] _GEN_12338 = 6'h23 == state ? $signed(temp) : $signed(_GEN_11826); // @[digest.scala 38:19 81:19]
  wire [31:0] _GEN_12339 = 6'h23 == state ? $signed(t) : $signed(_GEN_11828); // @[digest.scala 35:16 81:19]
  wire  _GEN_12340 = 6'h23 == state ? 1'h0 : _GEN_11829; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_12343 = 6'h23 == state ? $signed(e) : $signed(_GEN_11832); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_12344 = 6'h23 == state ? $signed(d) : $signed(_GEN_11833); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_12345 = 6'h23 == state ? $signed(c) : $signed(_GEN_11834); // @[digest.scala 26:16 81:19]
  wire  _GEN_12346 = 6'h23 == state ? 1'h0 : _GEN_11835; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_12349 = 6'h23 == state ? $signed(b) : $signed(_GEN_11838); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_12350 = 6'h23 == state ? $signed(a) : $signed(_GEN_11839); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_12351 = 6'h23 == state ? $signed(j) : $signed(_GEN_11840); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_12352 = 6'h23 == state ? $signed(i) : $signed(_GEN_11841); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_12434 = 6'h23 == state ? $signed(digest_0) : $signed(_GEN_11923); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12435 = 6'h23 == state ? $signed(digest_1) : $signed(_GEN_11924); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12436 = 6'h23 == state ? $signed(digest_2) : $signed(_GEN_11925); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12437 = 6'h23 == state ? $signed(digest_3) : $signed(_GEN_11926); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12438 = 6'h23 == state ? $signed(digest_4) : $signed(_GEN_11927); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12439 = 6'h23 == state ? $signed(digest_5) : $signed(_GEN_11928); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12440 = 6'h23 == state ? $signed(digest_6) : $signed(_GEN_11929); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12441 = 6'h23 == state ? $signed(digest_7) : $signed(_GEN_11930); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12442 = 6'h23 == state ? $signed(digest_8) : $signed(_GEN_11931); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12443 = 6'h23 == state ? $signed(digest_9) : $signed(_GEN_11932); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12444 = 6'h23 == state ? $signed(digest_10) : $signed(_GEN_11933); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12445 = 6'h23 == state ? $signed(digest_11) : $signed(_GEN_11934); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12446 = 6'h23 == state ? $signed(digest_12) : $signed(_GEN_11935); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12447 = 6'h23 == state ? $signed(digest_13) : $signed(_GEN_11936); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12448 = 6'h23 == state ? $signed(digest_14) : $signed(_GEN_11937); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12449 = 6'h23 == state ? $signed(digest_15) : $signed(_GEN_11938); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12450 = 6'h23 == state ? $signed(digest_16) : $signed(_GEN_11939); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12451 = 6'h23 == state ? $signed(digest_17) : $signed(_GEN_11940); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12452 = 6'h23 == state ? $signed(digest_18) : $signed(_GEN_11941); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12453 = 6'h23 == state ? $signed(digest_19) : $signed(_GEN_11942); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12454 = 6'h23 == state ? $signed(digest_20) : $signed(_GEN_11943); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12455 = 6'h23 == state ? $signed(digest_21) : $signed(_GEN_11944); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12456 = 6'h23 == state ? $signed(digest_22) : $signed(_GEN_11945); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12457 = 6'h23 == state ? $signed(digest_23) : $signed(_GEN_11946); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12458 = 6'h23 == state ? $signed(digest_24) : $signed(_GEN_11947); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12459 = 6'h23 == state ? $signed(digest_25) : $signed(_GEN_11948); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12460 = 6'h23 == state ? $signed(digest_26) : $signed(_GEN_11949); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12461 = 6'h23 == state ? $signed(digest_27) : $signed(_GEN_11950); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12462 = 6'h23 == state ? $signed(digest_28) : $signed(_GEN_11951); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12463 = 6'h23 == state ? $signed(digest_29) : $signed(_GEN_11952); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12464 = 6'h23 == state ? $signed(digest_30) : $signed(_GEN_11953); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12465 = 6'h23 == state ? $signed(digest_31) : $signed(_GEN_11954); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12466 = 6'h23 == state ? $signed(digest_32) : $signed(_GEN_11955); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12467 = 6'h23 == state ? $signed(digest_33) : $signed(_GEN_11956); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12468 = 6'h23 == state ? $signed(digest_34) : $signed(_GEN_11957); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12469 = 6'h23 == state ? $signed(digest_35) : $signed(_GEN_11958); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12470 = 6'h23 == state ? $signed(digest_36) : $signed(_GEN_11959); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12471 = 6'h23 == state ? $signed(digest_37) : $signed(_GEN_11960); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12472 = 6'h23 == state ? $signed(digest_38) : $signed(_GEN_11961); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12473 = 6'h23 == state ? $signed(digest_39) : $signed(_GEN_11962); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12474 = 6'h23 == state ? $signed(digest_40) : $signed(_GEN_11963); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12475 = 6'h23 == state ? $signed(digest_41) : $signed(_GEN_11964); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12476 = 6'h23 == state ? $signed(digest_42) : $signed(_GEN_11965); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12477 = 6'h23 == state ? $signed(digest_43) : $signed(_GEN_11966); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12478 = 6'h23 == state ? $signed(digest_44) : $signed(_GEN_11967); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12479 = 6'h23 == state ? $signed(digest_45) : $signed(_GEN_11968); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12480 = 6'h23 == state ? $signed(digest_46) : $signed(_GEN_11969); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12481 = 6'h23 == state ? $signed(digest_47) : $signed(_GEN_11970); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12482 = 6'h23 == state ? $signed(digest_48) : $signed(_GEN_11971); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12483 = 6'h23 == state ? $signed(digest_49) : $signed(_GEN_11972); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12484 = 6'h23 == state ? $signed(digest_50) : $signed(_GEN_11973); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12485 = 6'h23 == state ? $signed(digest_51) : $signed(_GEN_11974); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12486 = 6'h23 == state ? $signed(digest_52) : $signed(_GEN_11975); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12487 = 6'h23 == state ? $signed(digest_53) : $signed(_GEN_11976); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12488 = 6'h23 == state ? $signed(digest_54) : $signed(_GEN_11977); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12489 = 6'h23 == state ? $signed(digest_55) : $signed(_GEN_11978); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12490 = 6'h23 == state ? $signed(digest_56) : $signed(_GEN_11979); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12491 = 6'h23 == state ? $signed(digest_57) : $signed(_GEN_11980); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12492 = 6'h23 == state ? $signed(digest_58) : $signed(_GEN_11981); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12493 = 6'h23 == state ? $signed(digest_59) : $signed(_GEN_11982); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12494 = 6'h23 == state ? $signed(digest_60) : $signed(_GEN_11983); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12495 = 6'h23 == state ? $signed(digest_61) : $signed(_GEN_11984); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12496 = 6'h23 == state ? $signed(digest_62) : $signed(_GEN_11985); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12497 = 6'h23 == state ? $signed(digest_63) : $signed(_GEN_11986); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12498 = 6'h23 == state ? $signed(digest_64) : $signed(_GEN_11987); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12499 = 6'h23 == state ? $signed(digest_65) : $signed(_GEN_11988); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12500 = 6'h23 == state ? $signed(digest_66) : $signed(_GEN_11989); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12501 = 6'h23 == state ? $signed(digest_67) : $signed(_GEN_11990); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12502 = 6'h23 == state ? $signed(digest_68) : $signed(_GEN_11991); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12503 = 6'h23 == state ? $signed(digest_69) : $signed(_GEN_11992); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12504 = 6'h23 == state ? $signed(digest_70) : $signed(_GEN_11993); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12505 = 6'h23 == state ? $signed(digest_71) : $signed(_GEN_11994); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12506 = 6'h23 == state ? $signed(digest_72) : $signed(_GEN_11995); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12507 = 6'h23 == state ? $signed(digest_73) : $signed(_GEN_11996); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12508 = 6'h23 == state ? $signed(digest_74) : $signed(_GEN_11997); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12509 = 6'h23 == state ? $signed(digest_75) : $signed(_GEN_11998); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12510 = 6'h23 == state ? $signed(digest_76) : $signed(_GEN_11999); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12511 = 6'h23 == state ? $signed(digest_77) : $signed(_GEN_12000); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12512 = 6'h23 == state ? $signed(digest_78) : $signed(_GEN_12001); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12513 = 6'h23 == state ? $signed(digest_79) : $signed(_GEN_12002); // @[digest.scala 81:19 53:21]
  wire  _GEN_12515 = 6'h23 == state ? 1'h0 : _GEN_12004; // @[digest.scala 81:19 58:25]
  wire  _GEN_12598 = 6'h23 == state ? 1'h0 : _GEN_12087; // @[digest.scala 81:19 63:25]
  wire  _GEN_12681 = 6'h23 == state ? 1'h0 : _GEN_12170; // @[digest.scala 81:19 68:25]
  wire  _GEN_12764 = 6'h23 == state ? 1'h0 : _GEN_12253; // @[digest.scala 81:19 73:25]
  wire  _GEN_12847 = 6'h23 == state ? 1'h0 : _GEN_12336; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_12848 = 6'h22 == state ? $signed(_temp_T_61) : $signed(_GEN_12338); // @[digest.scala 219:18 81:19]
  wire [5:0] _GEN_12849 = 6'h22 == state ? 6'h28 : _GEN_12337; // @[digest.scala 220:19 81:19]
  wire [31:0] _GEN_12850 = 6'h22 == state ? $signed(t) : $signed(_GEN_12339); // @[digest.scala 35:16 81:19]
  wire  _GEN_12851 = 6'h22 == state ? 1'h0 : _GEN_12340; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_12854 = 6'h22 == state ? $signed(e) : $signed(_GEN_12343); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_12855 = 6'h22 == state ? $signed(d) : $signed(_GEN_12344); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_12856 = 6'h22 == state ? $signed(c) : $signed(_GEN_12345); // @[digest.scala 26:16 81:19]
  wire  _GEN_12857 = 6'h22 == state ? 1'h0 : _GEN_12346; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_12860 = 6'h22 == state ? $signed(b) : $signed(_GEN_12349); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_12861 = 6'h22 == state ? $signed(a) : $signed(_GEN_12350); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_12862 = 6'h22 == state ? $signed(j) : $signed(_GEN_12351); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_12863 = 6'h22 == state ? $signed(i) : $signed(_GEN_12352); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_12945 = 6'h22 == state ? $signed(digest_0) : $signed(_GEN_12434); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12946 = 6'h22 == state ? $signed(digest_1) : $signed(_GEN_12435); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12947 = 6'h22 == state ? $signed(digest_2) : $signed(_GEN_12436); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12948 = 6'h22 == state ? $signed(digest_3) : $signed(_GEN_12437); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12949 = 6'h22 == state ? $signed(digest_4) : $signed(_GEN_12438); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12950 = 6'h22 == state ? $signed(digest_5) : $signed(_GEN_12439); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12951 = 6'h22 == state ? $signed(digest_6) : $signed(_GEN_12440); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12952 = 6'h22 == state ? $signed(digest_7) : $signed(_GEN_12441); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12953 = 6'h22 == state ? $signed(digest_8) : $signed(_GEN_12442); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12954 = 6'h22 == state ? $signed(digest_9) : $signed(_GEN_12443); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12955 = 6'h22 == state ? $signed(digest_10) : $signed(_GEN_12444); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12956 = 6'h22 == state ? $signed(digest_11) : $signed(_GEN_12445); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12957 = 6'h22 == state ? $signed(digest_12) : $signed(_GEN_12446); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12958 = 6'h22 == state ? $signed(digest_13) : $signed(_GEN_12447); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12959 = 6'h22 == state ? $signed(digest_14) : $signed(_GEN_12448); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12960 = 6'h22 == state ? $signed(digest_15) : $signed(_GEN_12449); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12961 = 6'h22 == state ? $signed(digest_16) : $signed(_GEN_12450); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12962 = 6'h22 == state ? $signed(digest_17) : $signed(_GEN_12451); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12963 = 6'h22 == state ? $signed(digest_18) : $signed(_GEN_12452); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12964 = 6'h22 == state ? $signed(digest_19) : $signed(_GEN_12453); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12965 = 6'h22 == state ? $signed(digest_20) : $signed(_GEN_12454); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12966 = 6'h22 == state ? $signed(digest_21) : $signed(_GEN_12455); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12967 = 6'h22 == state ? $signed(digest_22) : $signed(_GEN_12456); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12968 = 6'h22 == state ? $signed(digest_23) : $signed(_GEN_12457); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12969 = 6'h22 == state ? $signed(digest_24) : $signed(_GEN_12458); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12970 = 6'h22 == state ? $signed(digest_25) : $signed(_GEN_12459); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12971 = 6'h22 == state ? $signed(digest_26) : $signed(_GEN_12460); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12972 = 6'h22 == state ? $signed(digest_27) : $signed(_GEN_12461); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12973 = 6'h22 == state ? $signed(digest_28) : $signed(_GEN_12462); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12974 = 6'h22 == state ? $signed(digest_29) : $signed(_GEN_12463); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12975 = 6'h22 == state ? $signed(digest_30) : $signed(_GEN_12464); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12976 = 6'h22 == state ? $signed(digest_31) : $signed(_GEN_12465); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12977 = 6'h22 == state ? $signed(digest_32) : $signed(_GEN_12466); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12978 = 6'h22 == state ? $signed(digest_33) : $signed(_GEN_12467); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12979 = 6'h22 == state ? $signed(digest_34) : $signed(_GEN_12468); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12980 = 6'h22 == state ? $signed(digest_35) : $signed(_GEN_12469); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12981 = 6'h22 == state ? $signed(digest_36) : $signed(_GEN_12470); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12982 = 6'h22 == state ? $signed(digest_37) : $signed(_GEN_12471); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12983 = 6'h22 == state ? $signed(digest_38) : $signed(_GEN_12472); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12984 = 6'h22 == state ? $signed(digest_39) : $signed(_GEN_12473); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12985 = 6'h22 == state ? $signed(digest_40) : $signed(_GEN_12474); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12986 = 6'h22 == state ? $signed(digest_41) : $signed(_GEN_12475); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12987 = 6'h22 == state ? $signed(digest_42) : $signed(_GEN_12476); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12988 = 6'h22 == state ? $signed(digest_43) : $signed(_GEN_12477); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12989 = 6'h22 == state ? $signed(digest_44) : $signed(_GEN_12478); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12990 = 6'h22 == state ? $signed(digest_45) : $signed(_GEN_12479); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12991 = 6'h22 == state ? $signed(digest_46) : $signed(_GEN_12480); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12992 = 6'h22 == state ? $signed(digest_47) : $signed(_GEN_12481); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12993 = 6'h22 == state ? $signed(digest_48) : $signed(_GEN_12482); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12994 = 6'h22 == state ? $signed(digest_49) : $signed(_GEN_12483); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12995 = 6'h22 == state ? $signed(digest_50) : $signed(_GEN_12484); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12996 = 6'h22 == state ? $signed(digest_51) : $signed(_GEN_12485); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12997 = 6'h22 == state ? $signed(digest_52) : $signed(_GEN_12486); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12998 = 6'h22 == state ? $signed(digest_53) : $signed(_GEN_12487); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_12999 = 6'h22 == state ? $signed(digest_54) : $signed(_GEN_12488); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13000 = 6'h22 == state ? $signed(digest_55) : $signed(_GEN_12489); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13001 = 6'h22 == state ? $signed(digest_56) : $signed(_GEN_12490); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13002 = 6'h22 == state ? $signed(digest_57) : $signed(_GEN_12491); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13003 = 6'h22 == state ? $signed(digest_58) : $signed(_GEN_12492); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13004 = 6'h22 == state ? $signed(digest_59) : $signed(_GEN_12493); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13005 = 6'h22 == state ? $signed(digest_60) : $signed(_GEN_12494); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13006 = 6'h22 == state ? $signed(digest_61) : $signed(_GEN_12495); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13007 = 6'h22 == state ? $signed(digest_62) : $signed(_GEN_12496); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13008 = 6'h22 == state ? $signed(digest_63) : $signed(_GEN_12497); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13009 = 6'h22 == state ? $signed(digest_64) : $signed(_GEN_12498); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13010 = 6'h22 == state ? $signed(digest_65) : $signed(_GEN_12499); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13011 = 6'h22 == state ? $signed(digest_66) : $signed(_GEN_12500); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13012 = 6'h22 == state ? $signed(digest_67) : $signed(_GEN_12501); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13013 = 6'h22 == state ? $signed(digest_68) : $signed(_GEN_12502); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13014 = 6'h22 == state ? $signed(digest_69) : $signed(_GEN_12503); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13015 = 6'h22 == state ? $signed(digest_70) : $signed(_GEN_12504); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13016 = 6'h22 == state ? $signed(digest_71) : $signed(_GEN_12505); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13017 = 6'h22 == state ? $signed(digest_72) : $signed(_GEN_12506); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13018 = 6'h22 == state ? $signed(digest_73) : $signed(_GEN_12507); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13019 = 6'h22 == state ? $signed(digest_74) : $signed(_GEN_12508); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13020 = 6'h22 == state ? $signed(digest_75) : $signed(_GEN_12509); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13021 = 6'h22 == state ? $signed(digest_76) : $signed(_GEN_12510); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13022 = 6'h22 == state ? $signed(digest_77) : $signed(_GEN_12511); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13023 = 6'h22 == state ? $signed(digest_78) : $signed(_GEN_12512); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13024 = 6'h22 == state ? $signed(digest_79) : $signed(_GEN_12513); // @[digest.scala 81:19 53:21]
  wire  _GEN_13026 = 6'h22 == state ? 1'h0 : _GEN_12515; // @[digest.scala 81:19 58:25]
  wire  _GEN_13109 = 6'h22 == state ? 1'h0 : _GEN_12598; // @[digest.scala 81:19 63:25]
  wire  _GEN_13192 = 6'h22 == state ? 1'h0 : _GEN_12681; // @[digest.scala 81:19 68:25]
  wire  _GEN_13275 = 6'h22 == state ? 1'h0 : _GEN_12764; // @[digest.scala 81:19 73:25]
  wire  _GEN_13358 = 6'h22 == state ? 1'h0 : _GEN_12847; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_13359 = 6'h21 == state ? $signed(_temp_T_58) : $signed(_GEN_12848); // @[digest.scala 215:18 81:19]
  wire [5:0] _GEN_13360 = 6'h21 == state ? 6'h22 : _GEN_12849; // @[digest.scala 216:19 81:19]
  wire [31:0] _GEN_13361 = 6'h21 == state ? $signed(t) : $signed(_GEN_12850); // @[digest.scala 35:16 81:19]
  wire  _GEN_13362 = 6'h21 == state ? 1'h0 : _GEN_12851; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_13365 = 6'h21 == state ? $signed(e) : $signed(_GEN_12854); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_13366 = 6'h21 == state ? $signed(d) : $signed(_GEN_12855); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_13367 = 6'h21 == state ? $signed(c) : $signed(_GEN_12856); // @[digest.scala 26:16 81:19]
  wire  _GEN_13368 = 6'h21 == state ? 1'h0 : _GEN_12857; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_13371 = 6'h21 == state ? $signed(b) : $signed(_GEN_12860); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_13372 = 6'h21 == state ? $signed(a) : $signed(_GEN_12861); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_13373 = 6'h21 == state ? $signed(j) : $signed(_GEN_12862); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_13374 = 6'h21 == state ? $signed(i) : $signed(_GEN_12863); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_13456 = 6'h21 == state ? $signed(digest_0) : $signed(_GEN_12945); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13457 = 6'h21 == state ? $signed(digest_1) : $signed(_GEN_12946); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13458 = 6'h21 == state ? $signed(digest_2) : $signed(_GEN_12947); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13459 = 6'h21 == state ? $signed(digest_3) : $signed(_GEN_12948); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13460 = 6'h21 == state ? $signed(digest_4) : $signed(_GEN_12949); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13461 = 6'h21 == state ? $signed(digest_5) : $signed(_GEN_12950); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13462 = 6'h21 == state ? $signed(digest_6) : $signed(_GEN_12951); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13463 = 6'h21 == state ? $signed(digest_7) : $signed(_GEN_12952); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13464 = 6'h21 == state ? $signed(digest_8) : $signed(_GEN_12953); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13465 = 6'h21 == state ? $signed(digest_9) : $signed(_GEN_12954); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13466 = 6'h21 == state ? $signed(digest_10) : $signed(_GEN_12955); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13467 = 6'h21 == state ? $signed(digest_11) : $signed(_GEN_12956); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13468 = 6'h21 == state ? $signed(digest_12) : $signed(_GEN_12957); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13469 = 6'h21 == state ? $signed(digest_13) : $signed(_GEN_12958); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13470 = 6'h21 == state ? $signed(digest_14) : $signed(_GEN_12959); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13471 = 6'h21 == state ? $signed(digest_15) : $signed(_GEN_12960); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13472 = 6'h21 == state ? $signed(digest_16) : $signed(_GEN_12961); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13473 = 6'h21 == state ? $signed(digest_17) : $signed(_GEN_12962); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13474 = 6'h21 == state ? $signed(digest_18) : $signed(_GEN_12963); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13475 = 6'h21 == state ? $signed(digest_19) : $signed(_GEN_12964); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13476 = 6'h21 == state ? $signed(digest_20) : $signed(_GEN_12965); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13477 = 6'h21 == state ? $signed(digest_21) : $signed(_GEN_12966); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13478 = 6'h21 == state ? $signed(digest_22) : $signed(_GEN_12967); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13479 = 6'h21 == state ? $signed(digest_23) : $signed(_GEN_12968); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13480 = 6'h21 == state ? $signed(digest_24) : $signed(_GEN_12969); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13481 = 6'h21 == state ? $signed(digest_25) : $signed(_GEN_12970); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13482 = 6'h21 == state ? $signed(digest_26) : $signed(_GEN_12971); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13483 = 6'h21 == state ? $signed(digest_27) : $signed(_GEN_12972); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13484 = 6'h21 == state ? $signed(digest_28) : $signed(_GEN_12973); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13485 = 6'h21 == state ? $signed(digest_29) : $signed(_GEN_12974); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13486 = 6'h21 == state ? $signed(digest_30) : $signed(_GEN_12975); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13487 = 6'h21 == state ? $signed(digest_31) : $signed(_GEN_12976); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13488 = 6'h21 == state ? $signed(digest_32) : $signed(_GEN_12977); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13489 = 6'h21 == state ? $signed(digest_33) : $signed(_GEN_12978); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13490 = 6'h21 == state ? $signed(digest_34) : $signed(_GEN_12979); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13491 = 6'h21 == state ? $signed(digest_35) : $signed(_GEN_12980); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13492 = 6'h21 == state ? $signed(digest_36) : $signed(_GEN_12981); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13493 = 6'h21 == state ? $signed(digest_37) : $signed(_GEN_12982); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13494 = 6'h21 == state ? $signed(digest_38) : $signed(_GEN_12983); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13495 = 6'h21 == state ? $signed(digest_39) : $signed(_GEN_12984); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13496 = 6'h21 == state ? $signed(digest_40) : $signed(_GEN_12985); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13497 = 6'h21 == state ? $signed(digest_41) : $signed(_GEN_12986); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13498 = 6'h21 == state ? $signed(digest_42) : $signed(_GEN_12987); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13499 = 6'h21 == state ? $signed(digest_43) : $signed(_GEN_12988); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13500 = 6'h21 == state ? $signed(digest_44) : $signed(_GEN_12989); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13501 = 6'h21 == state ? $signed(digest_45) : $signed(_GEN_12990); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13502 = 6'h21 == state ? $signed(digest_46) : $signed(_GEN_12991); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13503 = 6'h21 == state ? $signed(digest_47) : $signed(_GEN_12992); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13504 = 6'h21 == state ? $signed(digest_48) : $signed(_GEN_12993); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13505 = 6'h21 == state ? $signed(digest_49) : $signed(_GEN_12994); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13506 = 6'h21 == state ? $signed(digest_50) : $signed(_GEN_12995); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13507 = 6'h21 == state ? $signed(digest_51) : $signed(_GEN_12996); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13508 = 6'h21 == state ? $signed(digest_52) : $signed(_GEN_12997); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13509 = 6'h21 == state ? $signed(digest_53) : $signed(_GEN_12998); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13510 = 6'h21 == state ? $signed(digest_54) : $signed(_GEN_12999); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13511 = 6'h21 == state ? $signed(digest_55) : $signed(_GEN_13000); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13512 = 6'h21 == state ? $signed(digest_56) : $signed(_GEN_13001); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13513 = 6'h21 == state ? $signed(digest_57) : $signed(_GEN_13002); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13514 = 6'h21 == state ? $signed(digest_58) : $signed(_GEN_13003); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13515 = 6'h21 == state ? $signed(digest_59) : $signed(_GEN_13004); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13516 = 6'h21 == state ? $signed(digest_60) : $signed(_GEN_13005); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13517 = 6'h21 == state ? $signed(digest_61) : $signed(_GEN_13006); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13518 = 6'h21 == state ? $signed(digest_62) : $signed(_GEN_13007); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13519 = 6'h21 == state ? $signed(digest_63) : $signed(_GEN_13008); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13520 = 6'h21 == state ? $signed(digest_64) : $signed(_GEN_13009); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13521 = 6'h21 == state ? $signed(digest_65) : $signed(_GEN_13010); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13522 = 6'h21 == state ? $signed(digest_66) : $signed(_GEN_13011); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13523 = 6'h21 == state ? $signed(digest_67) : $signed(_GEN_13012); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13524 = 6'h21 == state ? $signed(digest_68) : $signed(_GEN_13013); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13525 = 6'h21 == state ? $signed(digest_69) : $signed(_GEN_13014); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13526 = 6'h21 == state ? $signed(digest_70) : $signed(_GEN_13015); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13527 = 6'h21 == state ? $signed(digest_71) : $signed(_GEN_13016); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13528 = 6'h21 == state ? $signed(digest_72) : $signed(_GEN_13017); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13529 = 6'h21 == state ? $signed(digest_73) : $signed(_GEN_13018); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13530 = 6'h21 == state ? $signed(digest_74) : $signed(_GEN_13019); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13531 = 6'h21 == state ? $signed(digest_75) : $signed(_GEN_13020); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13532 = 6'h21 == state ? $signed(digest_76) : $signed(_GEN_13021); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13533 = 6'h21 == state ? $signed(digest_77) : $signed(_GEN_13022); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13534 = 6'h21 == state ? $signed(digest_78) : $signed(_GEN_13023); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13535 = 6'h21 == state ? $signed(digest_79) : $signed(_GEN_13024); // @[digest.scala 81:19 53:21]
  wire  _GEN_13537 = 6'h21 == state ? 1'h0 : _GEN_13026; // @[digest.scala 81:19 58:25]
  wire  _GEN_13620 = 6'h21 == state ? 1'h0 : _GEN_13109; // @[digest.scala 81:19 63:25]
  wire  _GEN_13703 = 6'h21 == state ? 1'h0 : _GEN_13192; // @[digest.scala 81:19 68:25]
  wire  _GEN_13786 = 6'h21 == state ? 1'h0 : _GEN_13275; // @[digest.scala 81:19 73:25]
  wire  _GEN_13869 = 6'h21 == state ? 1'h0 : _GEN_13358; // @[digest.scala 81:19 78:25]
  wire [5:0] _GEN_13870 = 6'h20 == state ? _state_T_13 : _GEN_13360; // @[digest.scala 212:19 81:19]
  wire [31:0] _GEN_13871 = 6'h20 == state ? $signed(temp) : $signed(_GEN_13359); // @[digest.scala 38:19 81:19]
  wire [31:0] _GEN_13872 = 6'h20 == state ? $signed(t) : $signed(_GEN_13361); // @[digest.scala 35:16 81:19]
  wire  _GEN_13873 = 6'h20 == state ? 1'h0 : _GEN_13362; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_13876 = 6'h20 == state ? $signed(e) : $signed(_GEN_13365); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_13877 = 6'h20 == state ? $signed(d) : $signed(_GEN_13366); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_13878 = 6'h20 == state ? $signed(c) : $signed(_GEN_13367); // @[digest.scala 26:16 81:19]
  wire  _GEN_13879 = 6'h20 == state ? 1'h0 : _GEN_13368; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_13882 = 6'h20 == state ? $signed(b) : $signed(_GEN_13371); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_13883 = 6'h20 == state ? $signed(a) : $signed(_GEN_13372); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_13884 = 6'h20 == state ? $signed(j) : $signed(_GEN_13373); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_13885 = 6'h20 == state ? $signed(i) : $signed(_GEN_13374); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_13967 = 6'h20 == state ? $signed(digest_0) : $signed(_GEN_13456); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13968 = 6'h20 == state ? $signed(digest_1) : $signed(_GEN_13457); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13969 = 6'h20 == state ? $signed(digest_2) : $signed(_GEN_13458); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13970 = 6'h20 == state ? $signed(digest_3) : $signed(_GEN_13459); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13971 = 6'h20 == state ? $signed(digest_4) : $signed(_GEN_13460); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13972 = 6'h20 == state ? $signed(digest_5) : $signed(_GEN_13461); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13973 = 6'h20 == state ? $signed(digest_6) : $signed(_GEN_13462); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13974 = 6'h20 == state ? $signed(digest_7) : $signed(_GEN_13463); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13975 = 6'h20 == state ? $signed(digest_8) : $signed(_GEN_13464); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13976 = 6'h20 == state ? $signed(digest_9) : $signed(_GEN_13465); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13977 = 6'h20 == state ? $signed(digest_10) : $signed(_GEN_13466); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13978 = 6'h20 == state ? $signed(digest_11) : $signed(_GEN_13467); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13979 = 6'h20 == state ? $signed(digest_12) : $signed(_GEN_13468); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13980 = 6'h20 == state ? $signed(digest_13) : $signed(_GEN_13469); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13981 = 6'h20 == state ? $signed(digest_14) : $signed(_GEN_13470); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13982 = 6'h20 == state ? $signed(digest_15) : $signed(_GEN_13471); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13983 = 6'h20 == state ? $signed(digest_16) : $signed(_GEN_13472); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13984 = 6'h20 == state ? $signed(digest_17) : $signed(_GEN_13473); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13985 = 6'h20 == state ? $signed(digest_18) : $signed(_GEN_13474); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13986 = 6'h20 == state ? $signed(digest_19) : $signed(_GEN_13475); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13987 = 6'h20 == state ? $signed(digest_20) : $signed(_GEN_13476); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13988 = 6'h20 == state ? $signed(digest_21) : $signed(_GEN_13477); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13989 = 6'h20 == state ? $signed(digest_22) : $signed(_GEN_13478); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13990 = 6'h20 == state ? $signed(digest_23) : $signed(_GEN_13479); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13991 = 6'h20 == state ? $signed(digest_24) : $signed(_GEN_13480); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13992 = 6'h20 == state ? $signed(digest_25) : $signed(_GEN_13481); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13993 = 6'h20 == state ? $signed(digest_26) : $signed(_GEN_13482); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13994 = 6'h20 == state ? $signed(digest_27) : $signed(_GEN_13483); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13995 = 6'h20 == state ? $signed(digest_28) : $signed(_GEN_13484); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13996 = 6'h20 == state ? $signed(digest_29) : $signed(_GEN_13485); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13997 = 6'h20 == state ? $signed(digest_30) : $signed(_GEN_13486); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13998 = 6'h20 == state ? $signed(digest_31) : $signed(_GEN_13487); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_13999 = 6'h20 == state ? $signed(digest_32) : $signed(_GEN_13488); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14000 = 6'h20 == state ? $signed(digest_33) : $signed(_GEN_13489); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14001 = 6'h20 == state ? $signed(digest_34) : $signed(_GEN_13490); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14002 = 6'h20 == state ? $signed(digest_35) : $signed(_GEN_13491); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14003 = 6'h20 == state ? $signed(digest_36) : $signed(_GEN_13492); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14004 = 6'h20 == state ? $signed(digest_37) : $signed(_GEN_13493); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14005 = 6'h20 == state ? $signed(digest_38) : $signed(_GEN_13494); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14006 = 6'h20 == state ? $signed(digest_39) : $signed(_GEN_13495); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14007 = 6'h20 == state ? $signed(digest_40) : $signed(_GEN_13496); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14008 = 6'h20 == state ? $signed(digest_41) : $signed(_GEN_13497); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14009 = 6'h20 == state ? $signed(digest_42) : $signed(_GEN_13498); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14010 = 6'h20 == state ? $signed(digest_43) : $signed(_GEN_13499); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14011 = 6'h20 == state ? $signed(digest_44) : $signed(_GEN_13500); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14012 = 6'h20 == state ? $signed(digest_45) : $signed(_GEN_13501); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14013 = 6'h20 == state ? $signed(digest_46) : $signed(_GEN_13502); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14014 = 6'h20 == state ? $signed(digest_47) : $signed(_GEN_13503); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14015 = 6'h20 == state ? $signed(digest_48) : $signed(_GEN_13504); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14016 = 6'h20 == state ? $signed(digest_49) : $signed(_GEN_13505); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14017 = 6'h20 == state ? $signed(digest_50) : $signed(_GEN_13506); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14018 = 6'h20 == state ? $signed(digest_51) : $signed(_GEN_13507); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14019 = 6'h20 == state ? $signed(digest_52) : $signed(_GEN_13508); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14020 = 6'h20 == state ? $signed(digest_53) : $signed(_GEN_13509); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14021 = 6'h20 == state ? $signed(digest_54) : $signed(_GEN_13510); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14022 = 6'h20 == state ? $signed(digest_55) : $signed(_GEN_13511); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14023 = 6'h20 == state ? $signed(digest_56) : $signed(_GEN_13512); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14024 = 6'h20 == state ? $signed(digest_57) : $signed(_GEN_13513); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14025 = 6'h20 == state ? $signed(digest_58) : $signed(_GEN_13514); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14026 = 6'h20 == state ? $signed(digest_59) : $signed(_GEN_13515); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14027 = 6'h20 == state ? $signed(digest_60) : $signed(_GEN_13516); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14028 = 6'h20 == state ? $signed(digest_61) : $signed(_GEN_13517); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14029 = 6'h20 == state ? $signed(digest_62) : $signed(_GEN_13518); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14030 = 6'h20 == state ? $signed(digest_63) : $signed(_GEN_13519); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14031 = 6'h20 == state ? $signed(digest_64) : $signed(_GEN_13520); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14032 = 6'h20 == state ? $signed(digest_65) : $signed(_GEN_13521); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14033 = 6'h20 == state ? $signed(digest_66) : $signed(_GEN_13522); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14034 = 6'h20 == state ? $signed(digest_67) : $signed(_GEN_13523); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14035 = 6'h20 == state ? $signed(digest_68) : $signed(_GEN_13524); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14036 = 6'h20 == state ? $signed(digest_69) : $signed(_GEN_13525); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14037 = 6'h20 == state ? $signed(digest_70) : $signed(_GEN_13526); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14038 = 6'h20 == state ? $signed(digest_71) : $signed(_GEN_13527); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14039 = 6'h20 == state ? $signed(digest_72) : $signed(_GEN_13528); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14040 = 6'h20 == state ? $signed(digest_73) : $signed(_GEN_13529); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14041 = 6'h20 == state ? $signed(digest_74) : $signed(_GEN_13530); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14042 = 6'h20 == state ? $signed(digest_75) : $signed(_GEN_13531); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14043 = 6'h20 == state ? $signed(digest_76) : $signed(_GEN_13532); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14044 = 6'h20 == state ? $signed(digest_77) : $signed(_GEN_13533); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14045 = 6'h20 == state ? $signed(digest_78) : $signed(_GEN_13534); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14046 = 6'h20 == state ? $signed(digest_79) : $signed(_GEN_13535); // @[digest.scala 81:19 53:21]
  wire  _GEN_14048 = 6'h20 == state ? 1'h0 : _GEN_13537; // @[digest.scala 81:19 58:25]
  wire  _GEN_14131 = 6'h20 == state ? 1'h0 : _GEN_13620; // @[digest.scala 81:19 63:25]
  wire  _GEN_14214 = 6'h20 == state ? 1'h0 : _GEN_13703; // @[digest.scala 81:19 68:25]
  wire  _GEN_14297 = 6'h20 == state ? 1'h0 : _GEN_13786; // @[digest.scala 81:19 73:25]
  wire  _GEN_14380 = 6'h20 == state ? 1'h0 : _GEN_13869; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_14381 = 6'h1f == state ? $signed(_temp_T_54) : $signed(_GEN_13871); // @[digest.scala 208:18 81:19]
  wire [5:0] _GEN_14382 = 6'h1f == state ? 6'h28 : _GEN_13870; // @[digest.scala 209:19 81:19]
  wire [31:0] _GEN_14383 = 6'h1f == state ? $signed(t) : $signed(_GEN_13872); // @[digest.scala 35:16 81:19]
  wire  _GEN_14384 = 6'h1f == state ? 1'h0 : _GEN_13873; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_14387 = 6'h1f == state ? $signed(e) : $signed(_GEN_13876); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_14388 = 6'h1f == state ? $signed(d) : $signed(_GEN_13877); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_14389 = 6'h1f == state ? $signed(c) : $signed(_GEN_13878); // @[digest.scala 26:16 81:19]
  wire  _GEN_14390 = 6'h1f == state ? 1'h0 : _GEN_13879; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_14393 = 6'h1f == state ? $signed(b) : $signed(_GEN_13882); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_14394 = 6'h1f == state ? $signed(a) : $signed(_GEN_13883); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_14395 = 6'h1f == state ? $signed(j) : $signed(_GEN_13884); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_14396 = 6'h1f == state ? $signed(i) : $signed(_GEN_13885); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_14478 = 6'h1f == state ? $signed(digest_0) : $signed(_GEN_13967); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14479 = 6'h1f == state ? $signed(digest_1) : $signed(_GEN_13968); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14480 = 6'h1f == state ? $signed(digest_2) : $signed(_GEN_13969); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14481 = 6'h1f == state ? $signed(digest_3) : $signed(_GEN_13970); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14482 = 6'h1f == state ? $signed(digest_4) : $signed(_GEN_13971); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14483 = 6'h1f == state ? $signed(digest_5) : $signed(_GEN_13972); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14484 = 6'h1f == state ? $signed(digest_6) : $signed(_GEN_13973); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14485 = 6'h1f == state ? $signed(digest_7) : $signed(_GEN_13974); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14486 = 6'h1f == state ? $signed(digest_8) : $signed(_GEN_13975); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14487 = 6'h1f == state ? $signed(digest_9) : $signed(_GEN_13976); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14488 = 6'h1f == state ? $signed(digest_10) : $signed(_GEN_13977); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14489 = 6'h1f == state ? $signed(digest_11) : $signed(_GEN_13978); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14490 = 6'h1f == state ? $signed(digest_12) : $signed(_GEN_13979); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14491 = 6'h1f == state ? $signed(digest_13) : $signed(_GEN_13980); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14492 = 6'h1f == state ? $signed(digest_14) : $signed(_GEN_13981); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14493 = 6'h1f == state ? $signed(digest_15) : $signed(_GEN_13982); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14494 = 6'h1f == state ? $signed(digest_16) : $signed(_GEN_13983); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14495 = 6'h1f == state ? $signed(digest_17) : $signed(_GEN_13984); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14496 = 6'h1f == state ? $signed(digest_18) : $signed(_GEN_13985); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14497 = 6'h1f == state ? $signed(digest_19) : $signed(_GEN_13986); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14498 = 6'h1f == state ? $signed(digest_20) : $signed(_GEN_13987); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14499 = 6'h1f == state ? $signed(digest_21) : $signed(_GEN_13988); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14500 = 6'h1f == state ? $signed(digest_22) : $signed(_GEN_13989); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14501 = 6'h1f == state ? $signed(digest_23) : $signed(_GEN_13990); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14502 = 6'h1f == state ? $signed(digest_24) : $signed(_GEN_13991); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14503 = 6'h1f == state ? $signed(digest_25) : $signed(_GEN_13992); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14504 = 6'h1f == state ? $signed(digest_26) : $signed(_GEN_13993); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14505 = 6'h1f == state ? $signed(digest_27) : $signed(_GEN_13994); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14506 = 6'h1f == state ? $signed(digest_28) : $signed(_GEN_13995); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14507 = 6'h1f == state ? $signed(digest_29) : $signed(_GEN_13996); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14508 = 6'h1f == state ? $signed(digest_30) : $signed(_GEN_13997); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14509 = 6'h1f == state ? $signed(digest_31) : $signed(_GEN_13998); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14510 = 6'h1f == state ? $signed(digest_32) : $signed(_GEN_13999); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14511 = 6'h1f == state ? $signed(digest_33) : $signed(_GEN_14000); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14512 = 6'h1f == state ? $signed(digest_34) : $signed(_GEN_14001); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14513 = 6'h1f == state ? $signed(digest_35) : $signed(_GEN_14002); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14514 = 6'h1f == state ? $signed(digest_36) : $signed(_GEN_14003); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14515 = 6'h1f == state ? $signed(digest_37) : $signed(_GEN_14004); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14516 = 6'h1f == state ? $signed(digest_38) : $signed(_GEN_14005); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14517 = 6'h1f == state ? $signed(digest_39) : $signed(_GEN_14006); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14518 = 6'h1f == state ? $signed(digest_40) : $signed(_GEN_14007); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14519 = 6'h1f == state ? $signed(digest_41) : $signed(_GEN_14008); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14520 = 6'h1f == state ? $signed(digest_42) : $signed(_GEN_14009); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14521 = 6'h1f == state ? $signed(digest_43) : $signed(_GEN_14010); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14522 = 6'h1f == state ? $signed(digest_44) : $signed(_GEN_14011); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14523 = 6'h1f == state ? $signed(digest_45) : $signed(_GEN_14012); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14524 = 6'h1f == state ? $signed(digest_46) : $signed(_GEN_14013); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14525 = 6'h1f == state ? $signed(digest_47) : $signed(_GEN_14014); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14526 = 6'h1f == state ? $signed(digest_48) : $signed(_GEN_14015); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14527 = 6'h1f == state ? $signed(digest_49) : $signed(_GEN_14016); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14528 = 6'h1f == state ? $signed(digest_50) : $signed(_GEN_14017); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14529 = 6'h1f == state ? $signed(digest_51) : $signed(_GEN_14018); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14530 = 6'h1f == state ? $signed(digest_52) : $signed(_GEN_14019); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14531 = 6'h1f == state ? $signed(digest_53) : $signed(_GEN_14020); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14532 = 6'h1f == state ? $signed(digest_54) : $signed(_GEN_14021); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14533 = 6'h1f == state ? $signed(digest_55) : $signed(_GEN_14022); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14534 = 6'h1f == state ? $signed(digest_56) : $signed(_GEN_14023); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14535 = 6'h1f == state ? $signed(digest_57) : $signed(_GEN_14024); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14536 = 6'h1f == state ? $signed(digest_58) : $signed(_GEN_14025); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14537 = 6'h1f == state ? $signed(digest_59) : $signed(_GEN_14026); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14538 = 6'h1f == state ? $signed(digest_60) : $signed(_GEN_14027); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14539 = 6'h1f == state ? $signed(digest_61) : $signed(_GEN_14028); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14540 = 6'h1f == state ? $signed(digest_62) : $signed(_GEN_14029); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14541 = 6'h1f == state ? $signed(digest_63) : $signed(_GEN_14030); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14542 = 6'h1f == state ? $signed(digest_64) : $signed(_GEN_14031); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14543 = 6'h1f == state ? $signed(digest_65) : $signed(_GEN_14032); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14544 = 6'h1f == state ? $signed(digest_66) : $signed(_GEN_14033); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14545 = 6'h1f == state ? $signed(digest_67) : $signed(_GEN_14034); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14546 = 6'h1f == state ? $signed(digest_68) : $signed(_GEN_14035); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14547 = 6'h1f == state ? $signed(digest_69) : $signed(_GEN_14036); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14548 = 6'h1f == state ? $signed(digest_70) : $signed(_GEN_14037); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14549 = 6'h1f == state ? $signed(digest_71) : $signed(_GEN_14038); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14550 = 6'h1f == state ? $signed(digest_72) : $signed(_GEN_14039); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14551 = 6'h1f == state ? $signed(digest_73) : $signed(_GEN_14040); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14552 = 6'h1f == state ? $signed(digest_74) : $signed(_GEN_14041); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14553 = 6'h1f == state ? $signed(digest_75) : $signed(_GEN_14042); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14554 = 6'h1f == state ? $signed(digest_76) : $signed(_GEN_14043); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14555 = 6'h1f == state ? $signed(digest_77) : $signed(_GEN_14044); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14556 = 6'h1f == state ? $signed(digest_78) : $signed(_GEN_14045); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14557 = 6'h1f == state ? $signed(digest_79) : $signed(_GEN_14046); // @[digest.scala 81:19 53:21]
  wire  _GEN_14559 = 6'h1f == state ? 1'h0 : _GEN_14048; // @[digest.scala 81:19 58:25]
  wire  _GEN_14642 = 6'h1f == state ? 1'h0 : _GEN_14131; // @[digest.scala 81:19 63:25]
  wire  _GEN_14725 = 6'h1f == state ? 1'h0 : _GEN_14214; // @[digest.scala 81:19 68:25]
  wire  _GEN_14808 = 6'h1f == state ? 1'h0 : _GEN_14297; // @[digest.scala 81:19 73:25]
  wire  _GEN_14891 = 6'h1f == state ? 1'h0 : _GEN_14380; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_14892 = 6'h1e == state ? $signed(_temp_T_51) : $signed(_GEN_14381); // @[digest.scala 204:18 81:19]
  wire [5:0] _GEN_14893 = 6'h1e == state ? 6'h1f : _GEN_14382; // @[digest.scala 205:19 81:19]
  wire [31:0] _GEN_14894 = 6'h1e == state ? $signed(t) : $signed(_GEN_14383); // @[digest.scala 35:16 81:19]
  wire  _GEN_14895 = 6'h1e == state ? 1'h0 : _GEN_14384; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_14898 = 6'h1e == state ? $signed(e) : $signed(_GEN_14387); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_14899 = 6'h1e == state ? $signed(d) : $signed(_GEN_14388); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_14900 = 6'h1e == state ? $signed(c) : $signed(_GEN_14389); // @[digest.scala 26:16 81:19]
  wire  _GEN_14901 = 6'h1e == state ? 1'h0 : _GEN_14390; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_14904 = 6'h1e == state ? $signed(b) : $signed(_GEN_14393); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_14905 = 6'h1e == state ? $signed(a) : $signed(_GEN_14394); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_14906 = 6'h1e == state ? $signed(j) : $signed(_GEN_14395); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_14907 = 6'h1e == state ? $signed(i) : $signed(_GEN_14396); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_14989 = 6'h1e == state ? $signed(digest_0) : $signed(_GEN_14478); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14990 = 6'h1e == state ? $signed(digest_1) : $signed(_GEN_14479); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14991 = 6'h1e == state ? $signed(digest_2) : $signed(_GEN_14480); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14992 = 6'h1e == state ? $signed(digest_3) : $signed(_GEN_14481); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14993 = 6'h1e == state ? $signed(digest_4) : $signed(_GEN_14482); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14994 = 6'h1e == state ? $signed(digest_5) : $signed(_GEN_14483); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14995 = 6'h1e == state ? $signed(digest_6) : $signed(_GEN_14484); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14996 = 6'h1e == state ? $signed(digest_7) : $signed(_GEN_14485); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14997 = 6'h1e == state ? $signed(digest_8) : $signed(_GEN_14486); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14998 = 6'h1e == state ? $signed(digest_9) : $signed(_GEN_14487); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_14999 = 6'h1e == state ? $signed(digest_10) : $signed(_GEN_14488); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15000 = 6'h1e == state ? $signed(digest_11) : $signed(_GEN_14489); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15001 = 6'h1e == state ? $signed(digest_12) : $signed(_GEN_14490); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15002 = 6'h1e == state ? $signed(digest_13) : $signed(_GEN_14491); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15003 = 6'h1e == state ? $signed(digest_14) : $signed(_GEN_14492); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15004 = 6'h1e == state ? $signed(digest_15) : $signed(_GEN_14493); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15005 = 6'h1e == state ? $signed(digest_16) : $signed(_GEN_14494); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15006 = 6'h1e == state ? $signed(digest_17) : $signed(_GEN_14495); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15007 = 6'h1e == state ? $signed(digest_18) : $signed(_GEN_14496); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15008 = 6'h1e == state ? $signed(digest_19) : $signed(_GEN_14497); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15009 = 6'h1e == state ? $signed(digest_20) : $signed(_GEN_14498); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15010 = 6'h1e == state ? $signed(digest_21) : $signed(_GEN_14499); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15011 = 6'h1e == state ? $signed(digest_22) : $signed(_GEN_14500); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15012 = 6'h1e == state ? $signed(digest_23) : $signed(_GEN_14501); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15013 = 6'h1e == state ? $signed(digest_24) : $signed(_GEN_14502); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15014 = 6'h1e == state ? $signed(digest_25) : $signed(_GEN_14503); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15015 = 6'h1e == state ? $signed(digest_26) : $signed(_GEN_14504); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15016 = 6'h1e == state ? $signed(digest_27) : $signed(_GEN_14505); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15017 = 6'h1e == state ? $signed(digest_28) : $signed(_GEN_14506); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15018 = 6'h1e == state ? $signed(digest_29) : $signed(_GEN_14507); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15019 = 6'h1e == state ? $signed(digest_30) : $signed(_GEN_14508); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15020 = 6'h1e == state ? $signed(digest_31) : $signed(_GEN_14509); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15021 = 6'h1e == state ? $signed(digest_32) : $signed(_GEN_14510); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15022 = 6'h1e == state ? $signed(digest_33) : $signed(_GEN_14511); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15023 = 6'h1e == state ? $signed(digest_34) : $signed(_GEN_14512); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15024 = 6'h1e == state ? $signed(digest_35) : $signed(_GEN_14513); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15025 = 6'h1e == state ? $signed(digest_36) : $signed(_GEN_14514); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15026 = 6'h1e == state ? $signed(digest_37) : $signed(_GEN_14515); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15027 = 6'h1e == state ? $signed(digest_38) : $signed(_GEN_14516); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15028 = 6'h1e == state ? $signed(digest_39) : $signed(_GEN_14517); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15029 = 6'h1e == state ? $signed(digest_40) : $signed(_GEN_14518); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15030 = 6'h1e == state ? $signed(digest_41) : $signed(_GEN_14519); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15031 = 6'h1e == state ? $signed(digest_42) : $signed(_GEN_14520); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15032 = 6'h1e == state ? $signed(digest_43) : $signed(_GEN_14521); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15033 = 6'h1e == state ? $signed(digest_44) : $signed(_GEN_14522); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15034 = 6'h1e == state ? $signed(digest_45) : $signed(_GEN_14523); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15035 = 6'h1e == state ? $signed(digest_46) : $signed(_GEN_14524); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15036 = 6'h1e == state ? $signed(digest_47) : $signed(_GEN_14525); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15037 = 6'h1e == state ? $signed(digest_48) : $signed(_GEN_14526); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15038 = 6'h1e == state ? $signed(digest_49) : $signed(_GEN_14527); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15039 = 6'h1e == state ? $signed(digest_50) : $signed(_GEN_14528); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15040 = 6'h1e == state ? $signed(digest_51) : $signed(_GEN_14529); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15041 = 6'h1e == state ? $signed(digest_52) : $signed(_GEN_14530); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15042 = 6'h1e == state ? $signed(digest_53) : $signed(_GEN_14531); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15043 = 6'h1e == state ? $signed(digest_54) : $signed(_GEN_14532); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15044 = 6'h1e == state ? $signed(digest_55) : $signed(_GEN_14533); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15045 = 6'h1e == state ? $signed(digest_56) : $signed(_GEN_14534); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15046 = 6'h1e == state ? $signed(digest_57) : $signed(_GEN_14535); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15047 = 6'h1e == state ? $signed(digest_58) : $signed(_GEN_14536); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15048 = 6'h1e == state ? $signed(digest_59) : $signed(_GEN_14537); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15049 = 6'h1e == state ? $signed(digest_60) : $signed(_GEN_14538); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15050 = 6'h1e == state ? $signed(digest_61) : $signed(_GEN_14539); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15051 = 6'h1e == state ? $signed(digest_62) : $signed(_GEN_14540); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15052 = 6'h1e == state ? $signed(digest_63) : $signed(_GEN_14541); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15053 = 6'h1e == state ? $signed(digest_64) : $signed(_GEN_14542); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15054 = 6'h1e == state ? $signed(digest_65) : $signed(_GEN_14543); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15055 = 6'h1e == state ? $signed(digest_66) : $signed(_GEN_14544); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15056 = 6'h1e == state ? $signed(digest_67) : $signed(_GEN_14545); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15057 = 6'h1e == state ? $signed(digest_68) : $signed(_GEN_14546); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15058 = 6'h1e == state ? $signed(digest_69) : $signed(_GEN_14547); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15059 = 6'h1e == state ? $signed(digest_70) : $signed(_GEN_14548); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15060 = 6'h1e == state ? $signed(digest_71) : $signed(_GEN_14549); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15061 = 6'h1e == state ? $signed(digest_72) : $signed(_GEN_14550); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15062 = 6'h1e == state ? $signed(digest_73) : $signed(_GEN_14551); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15063 = 6'h1e == state ? $signed(digest_74) : $signed(_GEN_14552); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15064 = 6'h1e == state ? $signed(digest_75) : $signed(_GEN_14553); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15065 = 6'h1e == state ? $signed(digest_76) : $signed(_GEN_14554); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15066 = 6'h1e == state ? $signed(digest_77) : $signed(_GEN_14555); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15067 = 6'h1e == state ? $signed(digest_78) : $signed(_GEN_14556); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15068 = 6'h1e == state ? $signed(digest_79) : $signed(_GEN_14557); // @[digest.scala 81:19 53:21]
  wire  _GEN_15070 = 6'h1e == state ? 1'h0 : _GEN_14559; // @[digest.scala 81:19 58:25]
  wire  _GEN_15153 = 6'h1e == state ? 1'h0 : _GEN_14642; // @[digest.scala 81:19 63:25]
  wire  _GEN_15236 = 6'h1e == state ? 1'h0 : _GEN_14725; // @[digest.scala 81:19 68:25]
  wire  _GEN_15319 = 6'h1e == state ? 1'h0 : _GEN_14808; // @[digest.scala 81:19 73:25]
  wire  _GEN_15402 = 6'h1e == state ? 1'h0 : _GEN_14891; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_15403 = 6'h1d == state ? $signed(_temp_T_45) : $signed(_GEN_14892); // @[digest.scala 200:18 81:19]
  wire [5:0] _GEN_15404 = 6'h1d == state ? 6'h1e : _GEN_14893; // @[digest.scala 201:19 81:19]
  wire [31:0] _GEN_15405 = 6'h1d == state ? $signed(t) : $signed(_GEN_14894); // @[digest.scala 35:16 81:19]
  wire  _GEN_15406 = 6'h1d == state ? 1'h0 : _GEN_14895; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_15409 = 6'h1d == state ? $signed(e) : $signed(_GEN_14898); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_15410 = 6'h1d == state ? $signed(d) : $signed(_GEN_14899); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_15411 = 6'h1d == state ? $signed(c) : $signed(_GEN_14900); // @[digest.scala 26:16 81:19]
  wire  _GEN_15412 = 6'h1d == state ? 1'h0 : _GEN_14901; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_15415 = 6'h1d == state ? $signed(b) : $signed(_GEN_14904); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_15416 = 6'h1d == state ? $signed(a) : $signed(_GEN_14905); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_15417 = 6'h1d == state ? $signed(j) : $signed(_GEN_14906); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_15418 = 6'h1d == state ? $signed(i) : $signed(_GEN_14907); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_15500 = 6'h1d == state ? $signed(digest_0) : $signed(_GEN_14989); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15501 = 6'h1d == state ? $signed(digest_1) : $signed(_GEN_14990); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15502 = 6'h1d == state ? $signed(digest_2) : $signed(_GEN_14991); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15503 = 6'h1d == state ? $signed(digest_3) : $signed(_GEN_14992); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15504 = 6'h1d == state ? $signed(digest_4) : $signed(_GEN_14993); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15505 = 6'h1d == state ? $signed(digest_5) : $signed(_GEN_14994); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15506 = 6'h1d == state ? $signed(digest_6) : $signed(_GEN_14995); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15507 = 6'h1d == state ? $signed(digest_7) : $signed(_GEN_14996); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15508 = 6'h1d == state ? $signed(digest_8) : $signed(_GEN_14997); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15509 = 6'h1d == state ? $signed(digest_9) : $signed(_GEN_14998); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15510 = 6'h1d == state ? $signed(digest_10) : $signed(_GEN_14999); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15511 = 6'h1d == state ? $signed(digest_11) : $signed(_GEN_15000); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15512 = 6'h1d == state ? $signed(digest_12) : $signed(_GEN_15001); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15513 = 6'h1d == state ? $signed(digest_13) : $signed(_GEN_15002); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15514 = 6'h1d == state ? $signed(digest_14) : $signed(_GEN_15003); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15515 = 6'h1d == state ? $signed(digest_15) : $signed(_GEN_15004); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15516 = 6'h1d == state ? $signed(digest_16) : $signed(_GEN_15005); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15517 = 6'h1d == state ? $signed(digest_17) : $signed(_GEN_15006); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15518 = 6'h1d == state ? $signed(digest_18) : $signed(_GEN_15007); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15519 = 6'h1d == state ? $signed(digest_19) : $signed(_GEN_15008); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15520 = 6'h1d == state ? $signed(digest_20) : $signed(_GEN_15009); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15521 = 6'h1d == state ? $signed(digest_21) : $signed(_GEN_15010); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15522 = 6'h1d == state ? $signed(digest_22) : $signed(_GEN_15011); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15523 = 6'h1d == state ? $signed(digest_23) : $signed(_GEN_15012); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15524 = 6'h1d == state ? $signed(digest_24) : $signed(_GEN_15013); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15525 = 6'h1d == state ? $signed(digest_25) : $signed(_GEN_15014); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15526 = 6'h1d == state ? $signed(digest_26) : $signed(_GEN_15015); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15527 = 6'h1d == state ? $signed(digest_27) : $signed(_GEN_15016); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15528 = 6'h1d == state ? $signed(digest_28) : $signed(_GEN_15017); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15529 = 6'h1d == state ? $signed(digest_29) : $signed(_GEN_15018); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15530 = 6'h1d == state ? $signed(digest_30) : $signed(_GEN_15019); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15531 = 6'h1d == state ? $signed(digest_31) : $signed(_GEN_15020); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15532 = 6'h1d == state ? $signed(digest_32) : $signed(_GEN_15021); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15533 = 6'h1d == state ? $signed(digest_33) : $signed(_GEN_15022); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15534 = 6'h1d == state ? $signed(digest_34) : $signed(_GEN_15023); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15535 = 6'h1d == state ? $signed(digest_35) : $signed(_GEN_15024); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15536 = 6'h1d == state ? $signed(digest_36) : $signed(_GEN_15025); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15537 = 6'h1d == state ? $signed(digest_37) : $signed(_GEN_15026); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15538 = 6'h1d == state ? $signed(digest_38) : $signed(_GEN_15027); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15539 = 6'h1d == state ? $signed(digest_39) : $signed(_GEN_15028); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15540 = 6'h1d == state ? $signed(digest_40) : $signed(_GEN_15029); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15541 = 6'h1d == state ? $signed(digest_41) : $signed(_GEN_15030); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15542 = 6'h1d == state ? $signed(digest_42) : $signed(_GEN_15031); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15543 = 6'h1d == state ? $signed(digest_43) : $signed(_GEN_15032); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15544 = 6'h1d == state ? $signed(digest_44) : $signed(_GEN_15033); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15545 = 6'h1d == state ? $signed(digest_45) : $signed(_GEN_15034); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15546 = 6'h1d == state ? $signed(digest_46) : $signed(_GEN_15035); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15547 = 6'h1d == state ? $signed(digest_47) : $signed(_GEN_15036); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15548 = 6'h1d == state ? $signed(digest_48) : $signed(_GEN_15037); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15549 = 6'h1d == state ? $signed(digest_49) : $signed(_GEN_15038); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15550 = 6'h1d == state ? $signed(digest_50) : $signed(_GEN_15039); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15551 = 6'h1d == state ? $signed(digest_51) : $signed(_GEN_15040); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15552 = 6'h1d == state ? $signed(digest_52) : $signed(_GEN_15041); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15553 = 6'h1d == state ? $signed(digest_53) : $signed(_GEN_15042); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15554 = 6'h1d == state ? $signed(digest_54) : $signed(_GEN_15043); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15555 = 6'h1d == state ? $signed(digest_55) : $signed(_GEN_15044); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15556 = 6'h1d == state ? $signed(digest_56) : $signed(_GEN_15045); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15557 = 6'h1d == state ? $signed(digest_57) : $signed(_GEN_15046); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15558 = 6'h1d == state ? $signed(digest_58) : $signed(_GEN_15047); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15559 = 6'h1d == state ? $signed(digest_59) : $signed(_GEN_15048); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15560 = 6'h1d == state ? $signed(digest_60) : $signed(_GEN_15049); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15561 = 6'h1d == state ? $signed(digest_61) : $signed(_GEN_15050); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15562 = 6'h1d == state ? $signed(digest_62) : $signed(_GEN_15051); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15563 = 6'h1d == state ? $signed(digest_63) : $signed(_GEN_15052); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15564 = 6'h1d == state ? $signed(digest_64) : $signed(_GEN_15053); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15565 = 6'h1d == state ? $signed(digest_65) : $signed(_GEN_15054); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15566 = 6'h1d == state ? $signed(digest_66) : $signed(_GEN_15055); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15567 = 6'h1d == state ? $signed(digest_67) : $signed(_GEN_15056); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15568 = 6'h1d == state ? $signed(digest_68) : $signed(_GEN_15057); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15569 = 6'h1d == state ? $signed(digest_69) : $signed(_GEN_15058); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15570 = 6'h1d == state ? $signed(digest_70) : $signed(_GEN_15059); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15571 = 6'h1d == state ? $signed(digest_71) : $signed(_GEN_15060); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15572 = 6'h1d == state ? $signed(digest_72) : $signed(_GEN_15061); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15573 = 6'h1d == state ? $signed(digest_73) : $signed(_GEN_15062); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15574 = 6'h1d == state ? $signed(digest_74) : $signed(_GEN_15063); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15575 = 6'h1d == state ? $signed(digest_75) : $signed(_GEN_15064); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15576 = 6'h1d == state ? $signed(digest_76) : $signed(_GEN_15065); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15577 = 6'h1d == state ? $signed(digest_77) : $signed(_GEN_15066); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15578 = 6'h1d == state ? $signed(digest_78) : $signed(_GEN_15067); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_15579 = 6'h1d == state ? $signed(digest_79) : $signed(_GEN_15068); // @[digest.scala 81:19 53:21]
  wire  _GEN_15581 = 6'h1d == state ? 1'h0 : _GEN_15070; // @[digest.scala 81:19 58:25]
  wire  _GEN_15664 = 6'h1d == state ? 1'h0 : _GEN_15153; // @[digest.scala 81:19 63:25]
  wire  _GEN_15747 = 6'h1d == state ? 1'h0 : _GEN_15236; // @[digest.scala 81:19 68:25]
  wire  _GEN_15830 = 6'h1d == state ? 1'h0 : _GEN_15319; // @[digest.scala 81:19 73:25]
  wire  _GEN_15913 = 6'h1d == state ? 1'h0 : _GEN_15402; // @[digest.scala 81:19 78:25]
  wire [5:0] _GEN_15914 = 6'h1c == state ? _state_T_11 : _GEN_15404; // @[digest.scala 197:19 81:19]
  wire [31:0] _GEN_15915 = 6'h1c == state ? $signed(temp) : $signed(_GEN_15403); // @[digest.scala 38:19 81:19]
  wire [31:0] _GEN_15916 = 6'h1c == state ? $signed(t) : $signed(_GEN_15405); // @[digest.scala 35:16 81:19]
  wire  _GEN_15917 = 6'h1c == state ? 1'h0 : _GEN_15406; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_15920 = 6'h1c == state ? $signed(e) : $signed(_GEN_15409); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_15921 = 6'h1c == state ? $signed(d) : $signed(_GEN_15410); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_15922 = 6'h1c == state ? $signed(c) : $signed(_GEN_15411); // @[digest.scala 26:16 81:19]
  wire  _GEN_15923 = 6'h1c == state ? 1'h0 : _GEN_15412; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_15926 = 6'h1c == state ? $signed(b) : $signed(_GEN_15415); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_15927 = 6'h1c == state ? $signed(a) : $signed(_GEN_15416); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_15928 = 6'h1c == state ? $signed(j) : $signed(_GEN_15417); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_15929 = 6'h1c == state ? $signed(i) : $signed(_GEN_15418); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_16011 = 6'h1c == state ? $signed(digest_0) : $signed(_GEN_15500); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16012 = 6'h1c == state ? $signed(digest_1) : $signed(_GEN_15501); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16013 = 6'h1c == state ? $signed(digest_2) : $signed(_GEN_15502); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16014 = 6'h1c == state ? $signed(digest_3) : $signed(_GEN_15503); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16015 = 6'h1c == state ? $signed(digest_4) : $signed(_GEN_15504); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16016 = 6'h1c == state ? $signed(digest_5) : $signed(_GEN_15505); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16017 = 6'h1c == state ? $signed(digest_6) : $signed(_GEN_15506); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16018 = 6'h1c == state ? $signed(digest_7) : $signed(_GEN_15507); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16019 = 6'h1c == state ? $signed(digest_8) : $signed(_GEN_15508); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16020 = 6'h1c == state ? $signed(digest_9) : $signed(_GEN_15509); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16021 = 6'h1c == state ? $signed(digest_10) : $signed(_GEN_15510); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16022 = 6'h1c == state ? $signed(digest_11) : $signed(_GEN_15511); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16023 = 6'h1c == state ? $signed(digest_12) : $signed(_GEN_15512); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16024 = 6'h1c == state ? $signed(digest_13) : $signed(_GEN_15513); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16025 = 6'h1c == state ? $signed(digest_14) : $signed(_GEN_15514); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16026 = 6'h1c == state ? $signed(digest_15) : $signed(_GEN_15515); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16027 = 6'h1c == state ? $signed(digest_16) : $signed(_GEN_15516); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16028 = 6'h1c == state ? $signed(digest_17) : $signed(_GEN_15517); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16029 = 6'h1c == state ? $signed(digest_18) : $signed(_GEN_15518); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16030 = 6'h1c == state ? $signed(digest_19) : $signed(_GEN_15519); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16031 = 6'h1c == state ? $signed(digest_20) : $signed(_GEN_15520); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16032 = 6'h1c == state ? $signed(digest_21) : $signed(_GEN_15521); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16033 = 6'h1c == state ? $signed(digest_22) : $signed(_GEN_15522); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16034 = 6'h1c == state ? $signed(digest_23) : $signed(_GEN_15523); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16035 = 6'h1c == state ? $signed(digest_24) : $signed(_GEN_15524); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16036 = 6'h1c == state ? $signed(digest_25) : $signed(_GEN_15525); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16037 = 6'h1c == state ? $signed(digest_26) : $signed(_GEN_15526); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16038 = 6'h1c == state ? $signed(digest_27) : $signed(_GEN_15527); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16039 = 6'h1c == state ? $signed(digest_28) : $signed(_GEN_15528); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16040 = 6'h1c == state ? $signed(digest_29) : $signed(_GEN_15529); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16041 = 6'h1c == state ? $signed(digest_30) : $signed(_GEN_15530); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16042 = 6'h1c == state ? $signed(digest_31) : $signed(_GEN_15531); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16043 = 6'h1c == state ? $signed(digest_32) : $signed(_GEN_15532); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16044 = 6'h1c == state ? $signed(digest_33) : $signed(_GEN_15533); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16045 = 6'h1c == state ? $signed(digest_34) : $signed(_GEN_15534); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16046 = 6'h1c == state ? $signed(digest_35) : $signed(_GEN_15535); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16047 = 6'h1c == state ? $signed(digest_36) : $signed(_GEN_15536); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16048 = 6'h1c == state ? $signed(digest_37) : $signed(_GEN_15537); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16049 = 6'h1c == state ? $signed(digest_38) : $signed(_GEN_15538); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16050 = 6'h1c == state ? $signed(digest_39) : $signed(_GEN_15539); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16051 = 6'h1c == state ? $signed(digest_40) : $signed(_GEN_15540); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16052 = 6'h1c == state ? $signed(digest_41) : $signed(_GEN_15541); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16053 = 6'h1c == state ? $signed(digest_42) : $signed(_GEN_15542); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16054 = 6'h1c == state ? $signed(digest_43) : $signed(_GEN_15543); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16055 = 6'h1c == state ? $signed(digest_44) : $signed(_GEN_15544); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16056 = 6'h1c == state ? $signed(digest_45) : $signed(_GEN_15545); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16057 = 6'h1c == state ? $signed(digest_46) : $signed(_GEN_15546); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16058 = 6'h1c == state ? $signed(digest_47) : $signed(_GEN_15547); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16059 = 6'h1c == state ? $signed(digest_48) : $signed(_GEN_15548); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16060 = 6'h1c == state ? $signed(digest_49) : $signed(_GEN_15549); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16061 = 6'h1c == state ? $signed(digest_50) : $signed(_GEN_15550); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16062 = 6'h1c == state ? $signed(digest_51) : $signed(_GEN_15551); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16063 = 6'h1c == state ? $signed(digest_52) : $signed(_GEN_15552); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16064 = 6'h1c == state ? $signed(digest_53) : $signed(_GEN_15553); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16065 = 6'h1c == state ? $signed(digest_54) : $signed(_GEN_15554); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16066 = 6'h1c == state ? $signed(digest_55) : $signed(_GEN_15555); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16067 = 6'h1c == state ? $signed(digest_56) : $signed(_GEN_15556); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16068 = 6'h1c == state ? $signed(digest_57) : $signed(_GEN_15557); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16069 = 6'h1c == state ? $signed(digest_58) : $signed(_GEN_15558); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16070 = 6'h1c == state ? $signed(digest_59) : $signed(_GEN_15559); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16071 = 6'h1c == state ? $signed(digest_60) : $signed(_GEN_15560); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16072 = 6'h1c == state ? $signed(digest_61) : $signed(_GEN_15561); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16073 = 6'h1c == state ? $signed(digest_62) : $signed(_GEN_15562); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16074 = 6'h1c == state ? $signed(digest_63) : $signed(_GEN_15563); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16075 = 6'h1c == state ? $signed(digest_64) : $signed(_GEN_15564); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16076 = 6'h1c == state ? $signed(digest_65) : $signed(_GEN_15565); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16077 = 6'h1c == state ? $signed(digest_66) : $signed(_GEN_15566); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16078 = 6'h1c == state ? $signed(digest_67) : $signed(_GEN_15567); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16079 = 6'h1c == state ? $signed(digest_68) : $signed(_GEN_15568); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16080 = 6'h1c == state ? $signed(digest_69) : $signed(_GEN_15569); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16081 = 6'h1c == state ? $signed(digest_70) : $signed(_GEN_15570); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16082 = 6'h1c == state ? $signed(digest_71) : $signed(_GEN_15571); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16083 = 6'h1c == state ? $signed(digest_72) : $signed(_GEN_15572); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16084 = 6'h1c == state ? $signed(digest_73) : $signed(_GEN_15573); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16085 = 6'h1c == state ? $signed(digest_74) : $signed(_GEN_15574); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16086 = 6'h1c == state ? $signed(digest_75) : $signed(_GEN_15575); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16087 = 6'h1c == state ? $signed(digest_76) : $signed(_GEN_15576); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16088 = 6'h1c == state ? $signed(digest_77) : $signed(_GEN_15577); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16089 = 6'h1c == state ? $signed(digest_78) : $signed(_GEN_15578); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16090 = 6'h1c == state ? $signed(digest_79) : $signed(_GEN_15579); // @[digest.scala 81:19 53:21]
  wire  _GEN_16092 = 6'h1c == state ? 1'h0 : _GEN_15581; // @[digest.scala 81:19 58:25]
  wire  _GEN_16175 = 6'h1c == state ? 1'h0 : _GEN_15664; // @[digest.scala 81:19 63:25]
  wire  _GEN_16258 = 6'h1c == state ? 1'h0 : _GEN_15747; // @[digest.scala 81:19 68:25]
  wire  _GEN_16341 = 6'h1c == state ? 1'h0 : _GEN_15830; // @[digest.scala 81:19 73:25]
  wire  _GEN_16424 = 6'h1c == state ? 1'h0 : _GEN_15913; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_16425 = 6'h1b == state ? $signed(_GEN_1041) : $signed(w_0); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16426 = 6'h1b == state ? $signed(_GEN_1042) : $signed(w_1); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16427 = 6'h1b == state ? $signed(_GEN_1043) : $signed(w_2); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16428 = 6'h1b == state ? $signed(_GEN_1044) : $signed(w_3); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16429 = 6'h1b == state ? $signed(_GEN_1045) : $signed(w_4); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16430 = 6'h1b == state ? $signed(_GEN_1046) : $signed(w_5); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16431 = 6'h1b == state ? $signed(_GEN_1047) : $signed(w_6); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16432 = 6'h1b == state ? $signed(_GEN_1048) : $signed(w_7); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16433 = 6'h1b == state ? $signed(_GEN_1049) : $signed(w_8); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16434 = 6'h1b == state ? $signed(_GEN_1050) : $signed(w_9); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16435 = 6'h1b == state ? $signed(_GEN_1051) : $signed(w_10); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16436 = 6'h1b == state ? $signed(_GEN_1052) : $signed(w_11); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16437 = 6'h1b == state ? $signed(_GEN_1053) : $signed(w_12); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16438 = 6'h1b == state ? $signed(_GEN_1054) : $signed(w_13); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16439 = 6'h1b == state ? $signed(_GEN_1055) : $signed(w_14); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16440 = 6'h1b == state ? $signed(_GEN_1056) : $signed(w_15); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16441 = 6'h1b == state ? $signed(_GEN_1057) : $signed(w_16); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16442 = 6'h1b == state ? $signed(_GEN_1058) : $signed(w_17); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16443 = 6'h1b == state ? $signed(_GEN_1059) : $signed(w_18); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16444 = 6'h1b == state ? $signed(_GEN_1060) : $signed(w_19); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16445 = 6'h1b == state ? $signed(_GEN_1061) : $signed(w_20); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16446 = 6'h1b == state ? $signed(_GEN_1062) : $signed(w_21); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16447 = 6'h1b == state ? $signed(_GEN_1063) : $signed(w_22); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16448 = 6'h1b == state ? $signed(_GEN_1064) : $signed(w_23); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16449 = 6'h1b == state ? $signed(_GEN_1065) : $signed(w_24); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16450 = 6'h1b == state ? $signed(_GEN_1066) : $signed(w_25); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16451 = 6'h1b == state ? $signed(_GEN_1067) : $signed(w_26); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16452 = 6'h1b == state ? $signed(_GEN_1068) : $signed(w_27); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16453 = 6'h1b == state ? $signed(_GEN_1069) : $signed(w_28); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16454 = 6'h1b == state ? $signed(_GEN_1070) : $signed(w_29); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16455 = 6'h1b == state ? $signed(_GEN_1071) : $signed(w_30); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16456 = 6'h1b == state ? $signed(_GEN_1072) : $signed(w_31); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16457 = 6'h1b == state ? $signed(_GEN_1073) : $signed(w_32); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16458 = 6'h1b == state ? $signed(_GEN_1074) : $signed(w_33); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16459 = 6'h1b == state ? $signed(_GEN_1075) : $signed(w_34); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16460 = 6'h1b == state ? $signed(_GEN_1076) : $signed(w_35); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16461 = 6'h1b == state ? $signed(_GEN_1077) : $signed(w_36); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16462 = 6'h1b == state ? $signed(_GEN_1078) : $signed(w_37); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16463 = 6'h1b == state ? $signed(_GEN_1079) : $signed(w_38); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16464 = 6'h1b == state ? $signed(_GEN_1080) : $signed(w_39); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16465 = 6'h1b == state ? $signed(_GEN_1081) : $signed(w_40); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16466 = 6'h1b == state ? $signed(_GEN_1082) : $signed(w_41); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16467 = 6'h1b == state ? $signed(_GEN_1083) : $signed(w_42); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16468 = 6'h1b == state ? $signed(_GEN_1084) : $signed(w_43); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16469 = 6'h1b == state ? $signed(_GEN_1085) : $signed(w_44); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16470 = 6'h1b == state ? $signed(_GEN_1086) : $signed(w_45); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16471 = 6'h1b == state ? $signed(_GEN_1087) : $signed(w_46); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16472 = 6'h1b == state ? $signed(_GEN_1088) : $signed(w_47); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16473 = 6'h1b == state ? $signed(_GEN_1089) : $signed(w_48); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16474 = 6'h1b == state ? $signed(_GEN_1090) : $signed(w_49); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16475 = 6'h1b == state ? $signed(_GEN_1091) : $signed(w_50); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16476 = 6'h1b == state ? $signed(_GEN_1092) : $signed(w_51); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16477 = 6'h1b == state ? $signed(_GEN_1093) : $signed(w_52); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16478 = 6'h1b == state ? $signed(_GEN_1094) : $signed(w_53); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16479 = 6'h1b == state ? $signed(_GEN_1095) : $signed(w_54); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16480 = 6'h1b == state ? $signed(_GEN_1096) : $signed(w_55); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16481 = 6'h1b == state ? $signed(_GEN_1097) : $signed(w_56); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16482 = 6'h1b == state ? $signed(_GEN_1098) : $signed(w_57); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16483 = 6'h1b == state ? $signed(_GEN_1099) : $signed(w_58); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16484 = 6'h1b == state ? $signed(_GEN_1100) : $signed(w_59); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16485 = 6'h1b == state ? $signed(_GEN_1101) : $signed(w_60); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16486 = 6'h1b == state ? $signed(_GEN_1102) : $signed(w_61); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16487 = 6'h1b == state ? $signed(_GEN_1103) : $signed(w_62); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16488 = 6'h1b == state ? $signed(_GEN_1104) : $signed(w_63); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16489 = 6'h1b == state ? $signed(_GEN_1105) : $signed(w_64); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16490 = 6'h1b == state ? $signed(_GEN_1106) : $signed(w_65); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16491 = 6'h1b == state ? $signed(_GEN_1107) : $signed(w_66); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16492 = 6'h1b == state ? $signed(_GEN_1108) : $signed(w_67); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16493 = 6'h1b == state ? $signed(_GEN_1109) : $signed(w_68); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16494 = 6'h1b == state ? $signed(_GEN_1110) : $signed(w_69); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16495 = 6'h1b == state ? $signed(_GEN_1111) : $signed(w_70); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16496 = 6'h1b == state ? $signed(_GEN_1112) : $signed(w_71); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16497 = 6'h1b == state ? $signed(_GEN_1113) : $signed(w_72); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16498 = 6'h1b == state ? $signed(_GEN_1114) : $signed(w_73); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16499 = 6'h1b == state ? $signed(_GEN_1115) : $signed(w_74); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16500 = 6'h1b == state ? $signed(_GEN_1116) : $signed(w_75); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16501 = 6'h1b == state ? $signed(_GEN_1117) : $signed(w_76); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16502 = 6'h1b == state ? $signed(_GEN_1118) : $signed(w_77); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16503 = 6'h1b == state ? $signed(_GEN_1119) : $signed(w_78); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_16504 = 6'h1b == state ? $signed(_GEN_1120) : $signed(w_79); // @[digest.scala 40:16 81:19]
  wire  _GEN_16505 = 6'h1b == state & __m_rol_0_io_valid_T; // @[digest.scala 81:19 191:32 44:24]
  wire [5:0] _GEN_16508 = 6'h1b == state ? _state_T_9 : _GEN_15914; // @[digest.scala 194:19 81:19]
  wire [31:0] _GEN_16509 = 6'h1b == state ? $signed(temp) : $signed(_GEN_15915); // @[digest.scala 38:19 81:19]
  wire [31:0] _GEN_16510 = 6'h1b == state ? $signed(t) : $signed(_GEN_15916); // @[digest.scala 35:16 81:19]
  wire  _GEN_16511 = 6'h1b == state ? 1'h0 : _GEN_15917; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_16514 = 6'h1b == state ? $signed(e) : $signed(_GEN_15920); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_16515 = 6'h1b == state ? $signed(d) : $signed(_GEN_15921); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_16516 = 6'h1b == state ? $signed(c) : $signed(_GEN_15922); // @[digest.scala 26:16 81:19]
  wire  _GEN_16517 = 6'h1b == state ? 1'h0 : _GEN_15923; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_16520 = 6'h1b == state ? $signed(b) : $signed(_GEN_15926); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_16521 = 6'h1b == state ? $signed(a) : $signed(_GEN_15927); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_16522 = 6'h1b == state ? $signed(j) : $signed(_GEN_15928); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_16523 = 6'h1b == state ? $signed(i) : $signed(_GEN_15929); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_16605 = 6'h1b == state ? $signed(digest_0) : $signed(_GEN_16011); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16606 = 6'h1b == state ? $signed(digest_1) : $signed(_GEN_16012); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16607 = 6'h1b == state ? $signed(digest_2) : $signed(_GEN_16013); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16608 = 6'h1b == state ? $signed(digest_3) : $signed(_GEN_16014); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16609 = 6'h1b == state ? $signed(digest_4) : $signed(_GEN_16015); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16610 = 6'h1b == state ? $signed(digest_5) : $signed(_GEN_16016); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16611 = 6'h1b == state ? $signed(digest_6) : $signed(_GEN_16017); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16612 = 6'h1b == state ? $signed(digest_7) : $signed(_GEN_16018); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16613 = 6'h1b == state ? $signed(digest_8) : $signed(_GEN_16019); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16614 = 6'h1b == state ? $signed(digest_9) : $signed(_GEN_16020); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16615 = 6'h1b == state ? $signed(digest_10) : $signed(_GEN_16021); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16616 = 6'h1b == state ? $signed(digest_11) : $signed(_GEN_16022); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16617 = 6'h1b == state ? $signed(digest_12) : $signed(_GEN_16023); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16618 = 6'h1b == state ? $signed(digest_13) : $signed(_GEN_16024); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16619 = 6'h1b == state ? $signed(digest_14) : $signed(_GEN_16025); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16620 = 6'h1b == state ? $signed(digest_15) : $signed(_GEN_16026); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16621 = 6'h1b == state ? $signed(digest_16) : $signed(_GEN_16027); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16622 = 6'h1b == state ? $signed(digest_17) : $signed(_GEN_16028); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16623 = 6'h1b == state ? $signed(digest_18) : $signed(_GEN_16029); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16624 = 6'h1b == state ? $signed(digest_19) : $signed(_GEN_16030); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16625 = 6'h1b == state ? $signed(digest_20) : $signed(_GEN_16031); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16626 = 6'h1b == state ? $signed(digest_21) : $signed(_GEN_16032); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16627 = 6'h1b == state ? $signed(digest_22) : $signed(_GEN_16033); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16628 = 6'h1b == state ? $signed(digest_23) : $signed(_GEN_16034); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16629 = 6'h1b == state ? $signed(digest_24) : $signed(_GEN_16035); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16630 = 6'h1b == state ? $signed(digest_25) : $signed(_GEN_16036); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16631 = 6'h1b == state ? $signed(digest_26) : $signed(_GEN_16037); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16632 = 6'h1b == state ? $signed(digest_27) : $signed(_GEN_16038); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16633 = 6'h1b == state ? $signed(digest_28) : $signed(_GEN_16039); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16634 = 6'h1b == state ? $signed(digest_29) : $signed(_GEN_16040); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16635 = 6'h1b == state ? $signed(digest_30) : $signed(_GEN_16041); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16636 = 6'h1b == state ? $signed(digest_31) : $signed(_GEN_16042); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16637 = 6'h1b == state ? $signed(digest_32) : $signed(_GEN_16043); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16638 = 6'h1b == state ? $signed(digest_33) : $signed(_GEN_16044); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16639 = 6'h1b == state ? $signed(digest_34) : $signed(_GEN_16045); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16640 = 6'h1b == state ? $signed(digest_35) : $signed(_GEN_16046); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16641 = 6'h1b == state ? $signed(digest_36) : $signed(_GEN_16047); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16642 = 6'h1b == state ? $signed(digest_37) : $signed(_GEN_16048); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16643 = 6'h1b == state ? $signed(digest_38) : $signed(_GEN_16049); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16644 = 6'h1b == state ? $signed(digest_39) : $signed(_GEN_16050); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16645 = 6'h1b == state ? $signed(digest_40) : $signed(_GEN_16051); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16646 = 6'h1b == state ? $signed(digest_41) : $signed(_GEN_16052); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16647 = 6'h1b == state ? $signed(digest_42) : $signed(_GEN_16053); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16648 = 6'h1b == state ? $signed(digest_43) : $signed(_GEN_16054); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16649 = 6'h1b == state ? $signed(digest_44) : $signed(_GEN_16055); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16650 = 6'h1b == state ? $signed(digest_45) : $signed(_GEN_16056); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16651 = 6'h1b == state ? $signed(digest_46) : $signed(_GEN_16057); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16652 = 6'h1b == state ? $signed(digest_47) : $signed(_GEN_16058); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16653 = 6'h1b == state ? $signed(digest_48) : $signed(_GEN_16059); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16654 = 6'h1b == state ? $signed(digest_49) : $signed(_GEN_16060); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16655 = 6'h1b == state ? $signed(digest_50) : $signed(_GEN_16061); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16656 = 6'h1b == state ? $signed(digest_51) : $signed(_GEN_16062); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16657 = 6'h1b == state ? $signed(digest_52) : $signed(_GEN_16063); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16658 = 6'h1b == state ? $signed(digest_53) : $signed(_GEN_16064); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16659 = 6'h1b == state ? $signed(digest_54) : $signed(_GEN_16065); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16660 = 6'h1b == state ? $signed(digest_55) : $signed(_GEN_16066); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16661 = 6'h1b == state ? $signed(digest_56) : $signed(_GEN_16067); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16662 = 6'h1b == state ? $signed(digest_57) : $signed(_GEN_16068); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16663 = 6'h1b == state ? $signed(digest_58) : $signed(_GEN_16069); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16664 = 6'h1b == state ? $signed(digest_59) : $signed(_GEN_16070); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16665 = 6'h1b == state ? $signed(digest_60) : $signed(_GEN_16071); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16666 = 6'h1b == state ? $signed(digest_61) : $signed(_GEN_16072); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16667 = 6'h1b == state ? $signed(digest_62) : $signed(_GEN_16073); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16668 = 6'h1b == state ? $signed(digest_63) : $signed(_GEN_16074); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16669 = 6'h1b == state ? $signed(digest_64) : $signed(_GEN_16075); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16670 = 6'h1b == state ? $signed(digest_65) : $signed(_GEN_16076); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16671 = 6'h1b == state ? $signed(digest_66) : $signed(_GEN_16077); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16672 = 6'h1b == state ? $signed(digest_67) : $signed(_GEN_16078); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16673 = 6'h1b == state ? $signed(digest_68) : $signed(_GEN_16079); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16674 = 6'h1b == state ? $signed(digest_69) : $signed(_GEN_16080); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16675 = 6'h1b == state ? $signed(digest_70) : $signed(_GEN_16081); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16676 = 6'h1b == state ? $signed(digest_71) : $signed(_GEN_16082); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16677 = 6'h1b == state ? $signed(digest_72) : $signed(_GEN_16083); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16678 = 6'h1b == state ? $signed(digest_73) : $signed(_GEN_16084); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16679 = 6'h1b == state ? $signed(digest_74) : $signed(_GEN_16085); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16680 = 6'h1b == state ? $signed(digest_75) : $signed(_GEN_16086); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16681 = 6'h1b == state ? $signed(digest_76) : $signed(_GEN_16087); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16682 = 6'h1b == state ? $signed(digest_77) : $signed(_GEN_16088); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16683 = 6'h1b == state ? $signed(digest_78) : $signed(_GEN_16089); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_16684 = 6'h1b == state ? $signed(digest_79) : $signed(_GEN_16090); // @[digest.scala 81:19 53:21]
  wire  _GEN_16686 = 6'h1b == state ? 1'h0 : _GEN_16092; // @[digest.scala 81:19 58:25]
  wire  _GEN_16769 = 6'h1b == state ? 1'h0 : _GEN_16175; // @[digest.scala 81:19 63:25]
  wire  _GEN_16852 = 6'h1b == state ? 1'h0 : _GEN_16258; // @[digest.scala 81:19 68:25]
  wire  _GEN_16935 = 6'h1b == state ? 1'h0 : _GEN_16341; // @[digest.scala 81:19 73:25]
  wire  _GEN_17018 = 6'h1b == state ? 1'h0 : _GEN_16424; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_17019 = 6'h1a == state ? $signed(_temp_T_43) : $signed(_GEN_16509); // @[digest.scala 186:18 81:19]
  wire [5:0] _GEN_17020 = 6'h1a == state ? 6'h1b : _GEN_16508; // @[digest.scala 187:19 81:19]
  wire [31:0] _GEN_17021 = 6'h1a == state ? $signed(w_0) : $signed(_GEN_16425); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17022 = 6'h1a == state ? $signed(w_1) : $signed(_GEN_16426); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17023 = 6'h1a == state ? $signed(w_2) : $signed(_GEN_16427); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17024 = 6'h1a == state ? $signed(w_3) : $signed(_GEN_16428); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17025 = 6'h1a == state ? $signed(w_4) : $signed(_GEN_16429); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17026 = 6'h1a == state ? $signed(w_5) : $signed(_GEN_16430); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17027 = 6'h1a == state ? $signed(w_6) : $signed(_GEN_16431); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17028 = 6'h1a == state ? $signed(w_7) : $signed(_GEN_16432); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17029 = 6'h1a == state ? $signed(w_8) : $signed(_GEN_16433); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17030 = 6'h1a == state ? $signed(w_9) : $signed(_GEN_16434); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17031 = 6'h1a == state ? $signed(w_10) : $signed(_GEN_16435); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17032 = 6'h1a == state ? $signed(w_11) : $signed(_GEN_16436); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17033 = 6'h1a == state ? $signed(w_12) : $signed(_GEN_16437); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17034 = 6'h1a == state ? $signed(w_13) : $signed(_GEN_16438); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17035 = 6'h1a == state ? $signed(w_14) : $signed(_GEN_16439); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17036 = 6'h1a == state ? $signed(w_15) : $signed(_GEN_16440); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17037 = 6'h1a == state ? $signed(w_16) : $signed(_GEN_16441); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17038 = 6'h1a == state ? $signed(w_17) : $signed(_GEN_16442); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17039 = 6'h1a == state ? $signed(w_18) : $signed(_GEN_16443); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17040 = 6'h1a == state ? $signed(w_19) : $signed(_GEN_16444); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17041 = 6'h1a == state ? $signed(w_20) : $signed(_GEN_16445); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17042 = 6'h1a == state ? $signed(w_21) : $signed(_GEN_16446); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17043 = 6'h1a == state ? $signed(w_22) : $signed(_GEN_16447); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17044 = 6'h1a == state ? $signed(w_23) : $signed(_GEN_16448); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17045 = 6'h1a == state ? $signed(w_24) : $signed(_GEN_16449); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17046 = 6'h1a == state ? $signed(w_25) : $signed(_GEN_16450); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17047 = 6'h1a == state ? $signed(w_26) : $signed(_GEN_16451); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17048 = 6'h1a == state ? $signed(w_27) : $signed(_GEN_16452); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17049 = 6'h1a == state ? $signed(w_28) : $signed(_GEN_16453); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17050 = 6'h1a == state ? $signed(w_29) : $signed(_GEN_16454); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17051 = 6'h1a == state ? $signed(w_30) : $signed(_GEN_16455); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17052 = 6'h1a == state ? $signed(w_31) : $signed(_GEN_16456); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17053 = 6'h1a == state ? $signed(w_32) : $signed(_GEN_16457); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17054 = 6'h1a == state ? $signed(w_33) : $signed(_GEN_16458); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17055 = 6'h1a == state ? $signed(w_34) : $signed(_GEN_16459); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17056 = 6'h1a == state ? $signed(w_35) : $signed(_GEN_16460); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17057 = 6'h1a == state ? $signed(w_36) : $signed(_GEN_16461); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17058 = 6'h1a == state ? $signed(w_37) : $signed(_GEN_16462); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17059 = 6'h1a == state ? $signed(w_38) : $signed(_GEN_16463); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17060 = 6'h1a == state ? $signed(w_39) : $signed(_GEN_16464); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17061 = 6'h1a == state ? $signed(w_40) : $signed(_GEN_16465); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17062 = 6'h1a == state ? $signed(w_41) : $signed(_GEN_16466); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17063 = 6'h1a == state ? $signed(w_42) : $signed(_GEN_16467); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17064 = 6'h1a == state ? $signed(w_43) : $signed(_GEN_16468); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17065 = 6'h1a == state ? $signed(w_44) : $signed(_GEN_16469); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17066 = 6'h1a == state ? $signed(w_45) : $signed(_GEN_16470); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17067 = 6'h1a == state ? $signed(w_46) : $signed(_GEN_16471); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17068 = 6'h1a == state ? $signed(w_47) : $signed(_GEN_16472); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17069 = 6'h1a == state ? $signed(w_48) : $signed(_GEN_16473); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17070 = 6'h1a == state ? $signed(w_49) : $signed(_GEN_16474); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17071 = 6'h1a == state ? $signed(w_50) : $signed(_GEN_16475); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17072 = 6'h1a == state ? $signed(w_51) : $signed(_GEN_16476); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17073 = 6'h1a == state ? $signed(w_52) : $signed(_GEN_16477); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17074 = 6'h1a == state ? $signed(w_53) : $signed(_GEN_16478); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17075 = 6'h1a == state ? $signed(w_54) : $signed(_GEN_16479); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17076 = 6'h1a == state ? $signed(w_55) : $signed(_GEN_16480); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17077 = 6'h1a == state ? $signed(w_56) : $signed(_GEN_16481); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17078 = 6'h1a == state ? $signed(w_57) : $signed(_GEN_16482); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17079 = 6'h1a == state ? $signed(w_58) : $signed(_GEN_16483); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17080 = 6'h1a == state ? $signed(w_59) : $signed(_GEN_16484); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17081 = 6'h1a == state ? $signed(w_60) : $signed(_GEN_16485); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17082 = 6'h1a == state ? $signed(w_61) : $signed(_GEN_16486); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17083 = 6'h1a == state ? $signed(w_62) : $signed(_GEN_16487); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17084 = 6'h1a == state ? $signed(w_63) : $signed(_GEN_16488); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17085 = 6'h1a == state ? $signed(w_64) : $signed(_GEN_16489); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17086 = 6'h1a == state ? $signed(w_65) : $signed(_GEN_16490); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17087 = 6'h1a == state ? $signed(w_66) : $signed(_GEN_16491); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17088 = 6'h1a == state ? $signed(w_67) : $signed(_GEN_16492); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17089 = 6'h1a == state ? $signed(w_68) : $signed(_GEN_16493); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17090 = 6'h1a == state ? $signed(w_69) : $signed(_GEN_16494); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17091 = 6'h1a == state ? $signed(w_70) : $signed(_GEN_16495); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17092 = 6'h1a == state ? $signed(w_71) : $signed(_GEN_16496); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17093 = 6'h1a == state ? $signed(w_72) : $signed(_GEN_16497); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17094 = 6'h1a == state ? $signed(w_73) : $signed(_GEN_16498); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17095 = 6'h1a == state ? $signed(w_74) : $signed(_GEN_16499); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17096 = 6'h1a == state ? $signed(w_75) : $signed(_GEN_16500); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17097 = 6'h1a == state ? $signed(w_76) : $signed(_GEN_16501); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17098 = 6'h1a == state ? $signed(w_77) : $signed(_GEN_16502); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17099 = 6'h1a == state ? $signed(w_78) : $signed(_GEN_16503); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_17100 = 6'h1a == state ? $signed(w_79) : $signed(_GEN_16504); // @[digest.scala 40:16 81:19]
  wire  _GEN_17101 = 6'h1a == state ? 1'h0 : _GEN_16505; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_17104 = 6'h1a == state ? $signed(t) : $signed(_GEN_16510); // @[digest.scala 35:16 81:19]
  wire  _GEN_17105 = 6'h1a == state ? 1'h0 : _GEN_16511; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_17108 = 6'h1a == state ? $signed(e) : $signed(_GEN_16514); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_17109 = 6'h1a == state ? $signed(d) : $signed(_GEN_16515); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_17110 = 6'h1a == state ? $signed(c) : $signed(_GEN_16516); // @[digest.scala 26:16 81:19]
  wire  _GEN_17111 = 6'h1a == state ? 1'h0 : _GEN_16517; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_17114 = 6'h1a == state ? $signed(b) : $signed(_GEN_16520); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_17115 = 6'h1a == state ? $signed(a) : $signed(_GEN_16521); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_17116 = 6'h1a == state ? $signed(j) : $signed(_GEN_16522); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_17117 = 6'h1a == state ? $signed(i) : $signed(_GEN_16523); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_17199 = 6'h1a == state ? $signed(digest_0) : $signed(_GEN_16605); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17200 = 6'h1a == state ? $signed(digest_1) : $signed(_GEN_16606); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17201 = 6'h1a == state ? $signed(digest_2) : $signed(_GEN_16607); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17202 = 6'h1a == state ? $signed(digest_3) : $signed(_GEN_16608); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17203 = 6'h1a == state ? $signed(digest_4) : $signed(_GEN_16609); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17204 = 6'h1a == state ? $signed(digest_5) : $signed(_GEN_16610); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17205 = 6'h1a == state ? $signed(digest_6) : $signed(_GEN_16611); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17206 = 6'h1a == state ? $signed(digest_7) : $signed(_GEN_16612); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17207 = 6'h1a == state ? $signed(digest_8) : $signed(_GEN_16613); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17208 = 6'h1a == state ? $signed(digest_9) : $signed(_GEN_16614); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17209 = 6'h1a == state ? $signed(digest_10) : $signed(_GEN_16615); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17210 = 6'h1a == state ? $signed(digest_11) : $signed(_GEN_16616); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17211 = 6'h1a == state ? $signed(digest_12) : $signed(_GEN_16617); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17212 = 6'h1a == state ? $signed(digest_13) : $signed(_GEN_16618); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17213 = 6'h1a == state ? $signed(digest_14) : $signed(_GEN_16619); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17214 = 6'h1a == state ? $signed(digest_15) : $signed(_GEN_16620); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17215 = 6'h1a == state ? $signed(digest_16) : $signed(_GEN_16621); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17216 = 6'h1a == state ? $signed(digest_17) : $signed(_GEN_16622); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17217 = 6'h1a == state ? $signed(digest_18) : $signed(_GEN_16623); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17218 = 6'h1a == state ? $signed(digest_19) : $signed(_GEN_16624); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17219 = 6'h1a == state ? $signed(digest_20) : $signed(_GEN_16625); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17220 = 6'h1a == state ? $signed(digest_21) : $signed(_GEN_16626); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17221 = 6'h1a == state ? $signed(digest_22) : $signed(_GEN_16627); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17222 = 6'h1a == state ? $signed(digest_23) : $signed(_GEN_16628); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17223 = 6'h1a == state ? $signed(digest_24) : $signed(_GEN_16629); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17224 = 6'h1a == state ? $signed(digest_25) : $signed(_GEN_16630); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17225 = 6'h1a == state ? $signed(digest_26) : $signed(_GEN_16631); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17226 = 6'h1a == state ? $signed(digest_27) : $signed(_GEN_16632); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17227 = 6'h1a == state ? $signed(digest_28) : $signed(_GEN_16633); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17228 = 6'h1a == state ? $signed(digest_29) : $signed(_GEN_16634); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17229 = 6'h1a == state ? $signed(digest_30) : $signed(_GEN_16635); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17230 = 6'h1a == state ? $signed(digest_31) : $signed(_GEN_16636); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17231 = 6'h1a == state ? $signed(digest_32) : $signed(_GEN_16637); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17232 = 6'h1a == state ? $signed(digest_33) : $signed(_GEN_16638); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17233 = 6'h1a == state ? $signed(digest_34) : $signed(_GEN_16639); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17234 = 6'h1a == state ? $signed(digest_35) : $signed(_GEN_16640); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17235 = 6'h1a == state ? $signed(digest_36) : $signed(_GEN_16641); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17236 = 6'h1a == state ? $signed(digest_37) : $signed(_GEN_16642); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17237 = 6'h1a == state ? $signed(digest_38) : $signed(_GEN_16643); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17238 = 6'h1a == state ? $signed(digest_39) : $signed(_GEN_16644); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17239 = 6'h1a == state ? $signed(digest_40) : $signed(_GEN_16645); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17240 = 6'h1a == state ? $signed(digest_41) : $signed(_GEN_16646); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17241 = 6'h1a == state ? $signed(digest_42) : $signed(_GEN_16647); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17242 = 6'h1a == state ? $signed(digest_43) : $signed(_GEN_16648); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17243 = 6'h1a == state ? $signed(digest_44) : $signed(_GEN_16649); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17244 = 6'h1a == state ? $signed(digest_45) : $signed(_GEN_16650); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17245 = 6'h1a == state ? $signed(digest_46) : $signed(_GEN_16651); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17246 = 6'h1a == state ? $signed(digest_47) : $signed(_GEN_16652); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17247 = 6'h1a == state ? $signed(digest_48) : $signed(_GEN_16653); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17248 = 6'h1a == state ? $signed(digest_49) : $signed(_GEN_16654); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17249 = 6'h1a == state ? $signed(digest_50) : $signed(_GEN_16655); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17250 = 6'h1a == state ? $signed(digest_51) : $signed(_GEN_16656); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17251 = 6'h1a == state ? $signed(digest_52) : $signed(_GEN_16657); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17252 = 6'h1a == state ? $signed(digest_53) : $signed(_GEN_16658); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17253 = 6'h1a == state ? $signed(digest_54) : $signed(_GEN_16659); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17254 = 6'h1a == state ? $signed(digest_55) : $signed(_GEN_16660); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17255 = 6'h1a == state ? $signed(digest_56) : $signed(_GEN_16661); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17256 = 6'h1a == state ? $signed(digest_57) : $signed(_GEN_16662); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17257 = 6'h1a == state ? $signed(digest_58) : $signed(_GEN_16663); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17258 = 6'h1a == state ? $signed(digest_59) : $signed(_GEN_16664); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17259 = 6'h1a == state ? $signed(digest_60) : $signed(_GEN_16665); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17260 = 6'h1a == state ? $signed(digest_61) : $signed(_GEN_16666); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17261 = 6'h1a == state ? $signed(digest_62) : $signed(_GEN_16667); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17262 = 6'h1a == state ? $signed(digest_63) : $signed(_GEN_16668); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17263 = 6'h1a == state ? $signed(digest_64) : $signed(_GEN_16669); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17264 = 6'h1a == state ? $signed(digest_65) : $signed(_GEN_16670); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17265 = 6'h1a == state ? $signed(digest_66) : $signed(_GEN_16671); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17266 = 6'h1a == state ? $signed(digest_67) : $signed(_GEN_16672); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17267 = 6'h1a == state ? $signed(digest_68) : $signed(_GEN_16673); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17268 = 6'h1a == state ? $signed(digest_69) : $signed(_GEN_16674); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17269 = 6'h1a == state ? $signed(digest_70) : $signed(_GEN_16675); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17270 = 6'h1a == state ? $signed(digest_71) : $signed(_GEN_16676); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17271 = 6'h1a == state ? $signed(digest_72) : $signed(_GEN_16677); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17272 = 6'h1a == state ? $signed(digest_73) : $signed(_GEN_16678); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17273 = 6'h1a == state ? $signed(digest_74) : $signed(_GEN_16679); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17274 = 6'h1a == state ? $signed(digest_75) : $signed(_GEN_16680); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17275 = 6'h1a == state ? $signed(digest_76) : $signed(_GEN_16681); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17276 = 6'h1a == state ? $signed(digest_77) : $signed(_GEN_16682); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17277 = 6'h1a == state ? $signed(digest_78) : $signed(_GEN_16683); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17278 = 6'h1a == state ? $signed(digest_79) : $signed(_GEN_16684); // @[digest.scala 81:19 53:21]
  wire  _GEN_17280 = 6'h1a == state ? 1'h0 : _GEN_16686; // @[digest.scala 81:19 58:25]
  wire  _GEN_17363 = 6'h1a == state ? 1'h0 : _GEN_16769; // @[digest.scala 81:19 63:25]
  wire  _GEN_17446 = 6'h1a == state ? 1'h0 : _GEN_16852; // @[digest.scala 81:19 68:25]
  wire  _GEN_17529 = 6'h1a == state ? 1'h0 : _GEN_16935; // @[digest.scala 81:19 73:25]
  wire  _GEN_17612 = 6'h1a == state ? 1'h0 : _GEN_17018; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_17613 = 6'h19 == state ? $signed(_GEN_561) : $signed(_GEN_17021); // @[digest.scala 81:19]
  wire [31:0] _GEN_17614 = 6'h19 == state ? $signed(_GEN_562) : $signed(_GEN_17022); // @[digest.scala 81:19]
  wire [31:0] _GEN_17615 = 6'h19 == state ? $signed(_GEN_563) : $signed(_GEN_17023); // @[digest.scala 81:19]
  wire [31:0] _GEN_17616 = 6'h19 == state ? $signed(_GEN_564) : $signed(_GEN_17024); // @[digest.scala 81:19]
  wire [31:0] _GEN_17617 = 6'h19 == state ? $signed(_GEN_565) : $signed(_GEN_17025); // @[digest.scala 81:19]
  wire [31:0] _GEN_17618 = 6'h19 == state ? $signed(_GEN_566) : $signed(_GEN_17026); // @[digest.scala 81:19]
  wire [31:0] _GEN_17619 = 6'h19 == state ? $signed(_GEN_567) : $signed(_GEN_17027); // @[digest.scala 81:19]
  wire [31:0] _GEN_17620 = 6'h19 == state ? $signed(_GEN_568) : $signed(_GEN_17028); // @[digest.scala 81:19]
  wire [31:0] _GEN_17621 = 6'h19 == state ? $signed(_GEN_569) : $signed(_GEN_17029); // @[digest.scala 81:19]
  wire [31:0] _GEN_17622 = 6'h19 == state ? $signed(_GEN_570) : $signed(_GEN_17030); // @[digest.scala 81:19]
  wire [31:0] _GEN_17623 = 6'h19 == state ? $signed(_GEN_571) : $signed(_GEN_17031); // @[digest.scala 81:19]
  wire [31:0] _GEN_17624 = 6'h19 == state ? $signed(_GEN_572) : $signed(_GEN_17032); // @[digest.scala 81:19]
  wire [31:0] _GEN_17625 = 6'h19 == state ? $signed(_GEN_573) : $signed(_GEN_17033); // @[digest.scala 81:19]
  wire [31:0] _GEN_17626 = 6'h19 == state ? $signed(_GEN_574) : $signed(_GEN_17034); // @[digest.scala 81:19]
  wire [31:0] _GEN_17627 = 6'h19 == state ? $signed(_GEN_575) : $signed(_GEN_17035); // @[digest.scala 81:19]
  wire [31:0] _GEN_17628 = 6'h19 == state ? $signed(_GEN_576) : $signed(_GEN_17036); // @[digest.scala 81:19]
  wire [31:0] _GEN_17629 = 6'h19 == state ? $signed(_GEN_577) : $signed(_GEN_17037); // @[digest.scala 81:19]
  wire [31:0] _GEN_17630 = 6'h19 == state ? $signed(_GEN_578) : $signed(_GEN_17038); // @[digest.scala 81:19]
  wire [31:0] _GEN_17631 = 6'h19 == state ? $signed(_GEN_579) : $signed(_GEN_17039); // @[digest.scala 81:19]
  wire [31:0] _GEN_17632 = 6'h19 == state ? $signed(_GEN_580) : $signed(_GEN_17040); // @[digest.scala 81:19]
  wire [31:0] _GEN_17633 = 6'h19 == state ? $signed(_GEN_581) : $signed(_GEN_17041); // @[digest.scala 81:19]
  wire [31:0] _GEN_17634 = 6'h19 == state ? $signed(_GEN_582) : $signed(_GEN_17042); // @[digest.scala 81:19]
  wire [31:0] _GEN_17635 = 6'h19 == state ? $signed(_GEN_583) : $signed(_GEN_17043); // @[digest.scala 81:19]
  wire [31:0] _GEN_17636 = 6'h19 == state ? $signed(_GEN_584) : $signed(_GEN_17044); // @[digest.scala 81:19]
  wire [31:0] _GEN_17637 = 6'h19 == state ? $signed(_GEN_585) : $signed(_GEN_17045); // @[digest.scala 81:19]
  wire [31:0] _GEN_17638 = 6'h19 == state ? $signed(_GEN_586) : $signed(_GEN_17046); // @[digest.scala 81:19]
  wire [31:0] _GEN_17639 = 6'h19 == state ? $signed(_GEN_587) : $signed(_GEN_17047); // @[digest.scala 81:19]
  wire [31:0] _GEN_17640 = 6'h19 == state ? $signed(_GEN_588) : $signed(_GEN_17048); // @[digest.scala 81:19]
  wire [31:0] _GEN_17641 = 6'h19 == state ? $signed(_GEN_589) : $signed(_GEN_17049); // @[digest.scala 81:19]
  wire [31:0] _GEN_17642 = 6'h19 == state ? $signed(_GEN_590) : $signed(_GEN_17050); // @[digest.scala 81:19]
  wire [31:0] _GEN_17643 = 6'h19 == state ? $signed(_GEN_591) : $signed(_GEN_17051); // @[digest.scala 81:19]
  wire [31:0] _GEN_17644 = 6'h19 == state ? $signed(_GEN_592) : $signed(_GEN_17052); // @[digest.scala 81:19]
  wire [31:0] _GEN_17645 = 6'h19 == state ? $signed(_GEN_593) : $signed(_GEN_17053); // @[digest.scala 81:19]
  wire [31:0] _GEN_17646 = 6'h19 == state ? $signed(_GEN_594) : $signed(_GEN_17054); // @[digest.scala 81:19]
  wire [31:0] _GEN_17647 = 6'h19 == state ? $signed(_GEN_595) : $signed(_GEN_17055); // @[digest.scala 81:19]
  wire [31:0] _GEN_17648 = 6'h19 == state ? $signed(_GEN_596) : $signed(_GEN_17056); // @[digest.scala 81:19]
  wire [31:0] _GEN_17649 = 6'h19 == state ? $signed(_GEN_597) : $signed(_GEN_17057); // @[digest.scala 81:19]
  wire [31:0] _GEN_17650 = 6'h19 == state ? $signed(_GEN_598) : $signed(_GEN_17058); // @[digest.scala 81:19]
  wire [31:0] _GEN_17651 = 6'h19 == state ? $signed(_GEN_599) : $signed(_GEN_17059); // @[digest.scala 81:19]
  wire [31:0] _GEN_17652 = 6'h19 == state ? $signed(_GEN_600) : $signed(_GEN_17060); // @[digest.scala 81:19]
  wire [31:0] _GEN_17653 = 6'h19 == state ? $signed(_GEN_601) : $signed(_GEN_17061); // @[digest.scala 81:19]
  wire [31:0] _GEN_17654 = 6'h19 == state ? $signed(_GEN_602) : $signed(_GEN_17062); // @[digest.scala 81:19]
  wire [31:0] _GEN_17655 = 6'h19 == state ? $signed(_GEN_603) : $signed(_GEN_17063); // @[digest.scala 81:19]
  wire [31:0] _GEN_17656 = 6'h19 == state ? $signed(_GEN_604) : $signed(_GEN_17064); // @[digest.scala 81:19]
  wire [31:0] _GEN_17657 = 6'h19 == state ? $signed(_GEN_605) : $signed(_GEN_17065); // @[digest.scala 81:19]
  wire [31:0] _GEN_17658 = 6'h19 == state ? $signed(_GEN_606) : $signed(_GEN_17066); // @[digest.scala 81:19]
  wire [31:0] _GEN_17659 = 6'h19 == state ? $signed(_GEN_607) : $signed(_GEN_17067); // @[digest.scala 81:19]
  wire [31:0] _GEN_17660 = 6'h19 == state ? $signed(_GEN_608) : $signed(_GEN_17068); // @[digest.scala 81:19]
  wire [31:0] _GEN_17661 = 6'h19 == state ? $signed(_GEN_609) : $signed(_GEN_17069); // @[digest.scala 81:19]
  wire [31:0] _GEN_17662 = 6'h19 == state ? $signed(_GEN_610) : $signed(_GEN_17070); // @[digest.scala 81:19]
  wire [31:0] _GEN_17663 = 6'h19 == state ? $signed(_GEN_611) : $signed(_GEN_17071); // @[digest.scala 81:19]
  wire [31:0] _GEN_17664 = 6'h19 == state ? $signed(_GEN_612) : $signed(_GEN_17072); // @[digest.scala 81:19]
  wire [31:0] _GEN_17665 = 6'h19 == state ? $signed(_GEN_613) : $signed(_GEN_17073); // @[digest.scala 81:19]
  wire [31:0] _GEN_17666 = 6'h19 == state ? $signed(_GEN_614) : $signed(_GEN_17074); // @[digest.scala 81:19]
  wire [31:0] _GEN_17667 = 6'h19 == state ? $signed(_GEN_615) : $signed(_GEN_17075); // @[digest.scala 81:19]
  wire [31:0] _GEN_17668 = 6'h19 == state ? $signed(_GEN_616) : $signed(_GEN_17076); // @[digest.scala 81:19]
  wire [31:0] _GEN_17669 = 6'h19 == state ? $signed(_GEN_617) : $signed(_GEN_17077); // @[digest.scala 81:19]
  wire [31:0] _GEN_17670 = 6'h19 == state ? $signed(_GEN_618) : $signed(_GEN_17078); // @[digest.scala 81:19]
  wire [31:0] _GEN_17671 = 6'h19 == state ? $signed(_GEN_619) : $signed(_GEN_17079); // @[digest.scala 81:19]
  wire [31:0] _GEN_17672 = 6'h19 == state ? $signed(_GEN_620) : $signed(_GEN_17080); // @[digest.scala 81:19]
  wire [31:0] _GEN_17673 = 6'h19 == state ? $signed(_GEN_621) : $signed(_GEN_17081); // @[digest.scala 81:19]
  wire [31:0] _GEN_17674 = 6'h19 == state ? $signed(_GEN_622) : $signed(_GEN_17082); // @[digest.scala 81:19]
  wire [31:0] _GEN_17675 = 6'h19 == state ? $signed(_GEN_623) : $signed(_GEN_17083); // @[digest.scala 81:19]
  wire [31:0] _GEN_17676 = 6'h19 == state ? $signed(_GEN_624) : $signed(_GEN_17084); // @[digest.scala 81:19]
  wire [31:0] _GEN_17677 = 6'h19 == state ? $signed(_GEN_625) : $signed(_GEN_17085); // @[digest.scala 81:19]
  wire [31:0] _GEN_17678 = 6'h19 == state ? $signed(_GEN_626) : $signed(_GEN_17086); // @[digest.scala 81:19]
  wire [31:0] _GEN_17679 = 6'h19 == state ? $signed(_GEN_627) : $signed(_GEN_17087); // @[digest.scala 81:19]
  wire [31:0] _GEN_17680 = 6'h19 == state ? $signed(_GEN_628) : $signed(_GEN_17088); // @[digest.scala 81:19]
  wire [31:0] _GEN_17681 = 6'h19 == state ? $signed(_GEN_629) : $signed(_GEN_17089); // @[digest.scala 81:19]
  wire [31:0] _GEN_17682 = 6'h19 == state ? $signed(_GEN_630) : $signed(_GEN_17090); // @[digest.scala 81:19]
  wire [31:0] _GEN_17683 = 6'h19 == state ? $signed(_GEN_631) : $signed(_GEN_17091); // @[digest.scala 81:19]
  wire [31:0] _GEN_17684 = 6'h19 == state ? $signed(_GEN_632) : $signed(_GEN_17092); // @[digest.scala 81:19]
  wire [31:0] _GEN_17685 = 6'h19 == state ? $signed(_GEN_633) : $signed(_GEN_17093); // @[digest.scala 81:19]
  wire [31:0] _GEN_17686 = 6'h19 == state ? $signed(_GEN_634) : $signed(_GEN_17094); // @[digest.scala 81:19]
  wire [31:0] _GEN_17687 = 6'h19 == state ? $signed(_GEN_635) : $signed(_GEN_17095); // @[digest.scala 81:19]
  wire [31:0] _GEN_17688 = 6'h19 == state ? $signed(_GEN_636) : $signed(_GEN_17096); // @[digest.scala 81:19]
  wire [31:0] _GEN_17689 = 6'h19 == state ? $signed(_GEN_637) : $signed(_GEN_17097); // @[digest.scala 81:19]
  wire [31:0] _GEN_17690 = 6'h19 == state ? $signed(_GEN_638) : $signed(_GEN_17098); // @[digest.scala 81:19]
  wire [31:0] _GEN_17691 = 6'h19 == state ? $signed(_GEN_639) : $signed(_GEN_17099); // @[digest.scala 81:19]
  wire [31:0] _GEN_17692 = 6'h19 == state ? $signed(_GEN_640) : $signed(_GEN_17100); // @[digest.scala 81:19]
  wire [5:0] _GEN_17693 = 6'h19 == state ? 6'h1c : _GEN_17020; // @[digest.scala 183:19 81:19]
  wire [31:0] _GEN_17694 = 6'h19 == state ? $signed(temp) : $signed(_GEN_17019); // @[digest.scala 38:19 81:19]
  wire  _GEN_17695 = 6'h19 == state ? 1'h0 : _GEN_17101; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_17698 = 6'h19 == state ? $signed(t) : $signed(_GEN_17104); // @[digest.scala 35:16 81:19]
  wire  _GEN_17699 = 6'h19 == state ? 1'h0 : _GEN_17105; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_17702 = 6'h19 == state ? $signed(e) : $signed(_GEN_17108); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_17703 = 6'h19 == state ? $signed(d) : $signed(_GEN_17109); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_17704 = 6'h19 == state ? $signed(c) : $signed(_GEN_17110); // @[digest.scala 26:16 81:19]
  wire  _GEN_17705 = 6'h19 == state ? 1'h0 : _GEN_17111; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_17708 = 6'h19 == state ? $signed(b) : $signed(_GEN_17114); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_17709 = 6'h19 == state ? $signed(a) : $signed(_GEN_17115); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_17710 = 6'h19 == state ? $signed(j) : $signed(_GEN_17116); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_17711 = 6'h19 == state ? $signed(i) : $signed(_GEN_17117); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_17793 = 6'h19 == state ? $signed(digest_0) : $signed(_GEN_17199); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17794 = 6'h19 == state ? $signed(digest_1) : $signed(_GEN_17200); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17795 = 6'h19 == state ? $signed(digest_2) : $signed(_GEN_17201); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17796 = 6'h19 == state ? $signed(digest_3) : $signed(_GEN_17202); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17797 = 6'h19 == state ? $signed(digest_4) : $signed(_GEN_17203); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17798 = 6'h19 == state ? $signed(digest_5) : $signed(_GEN_17204); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17799 = 6'h19 == state ? $signed(digest_6) : $signed(_GEN_17205); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17800 = 6'h19 == state ? $signed(digest_7) : $signed(_GEN_17206); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17801 = 6'h19 == state ? $signed(digest_8) : $signed(_GEN_17207); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17802 = 6'h19 == state ? $signed(digest_9) : $signed(_GEN_17208); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17803 = 6'h19 == state ? $signed(digest_10) : $signed(_GEN_17209); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17804 = 6'h19 == state ? $signed(digest_11) : $signed(_GEN_17210); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17805 = 6'h19 == state ? $signed(digest_12) : $signed(_GEN_17211); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17806 = 6'h19 == state ? $signed(digest_13) : $signed(_GEN_17212); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17807 = 6'h19 == state ? $signed(digest_14) : $signed(_GEN_17213); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17808 = 6'h19 == state ? $signed(digest_15) : $signed(_GEN_17214); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17809 = 6'h19 == state ? $signed(digest_16) : $signed(_GEN_17215); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17810 = 6'h19 == state ? $signed(digest_17) : $signed(_GEN_17216); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17811 = 6'h19 == state ? $signed(digest_18) : $signed(_GEN_17217); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17812 = 6'h19 == state ? $signed(digest_19) : $signed(_GEN_17218); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17813 = 6'h19 == state ? $signed(digest_20) : $signed(_GEN_17219); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17814 = 6'h19 == state ? $signed(digest_21) : $signed(_GEN_17220); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17815 = 6'h19 == state ? $signed(digest_22) : $signed(_GEN_17221); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17816 = 6'h19 == state ? $signed(digest_23) : $signed(_GEN_17222); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17817 = 6'h19 == state ? $signed(digest_24) : $signed(_GEN_17223); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17818 = 6'h19 == state ? $signed(digest_25) : $signed(_GEN_17224); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17819 = 6'h19 == state ? $signed(digest_26) : $signed(_GEN_17225); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17820 = 6'h19 == state ? $signed(digest_27) : $signed(_GEN_17226); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17821 = 6'h19 == state ? $signed(digest_28) : $signed(_GEN_17227); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17822 = 6'h19 == state ? $signed(digest_29) : $signed(_GEN_17228); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17823 = 6'h19 == state ? $signed(digest_30) : $signed(_GEN_17229); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17824 = 6'h19 == state ? $signed(digest_31) : $signed(_GEN_17230); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17825 = 6'h19 == state ? $signed(digest_32) : $signed(_GEN_17231); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17826 = 6'h19 == state ? $signed(digest_33) : $signed(_GEN_17232); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17827 = 6'h19 == state ? $signed(digest_34) : $signed(_GEN_17233); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17828 = 6'h19 == state ? $signed(digest_35) : $signed(_GEN_17234); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17829 = 6'h19 == state ? $signed(digest_36) : $signed(_GEN_17235); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17830 = 6'h19 == state ? $signed(digest_37) : $signed(_GEN_17236); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17831 = 6'h19 == state ? $signed(digest_38) : $signed(_GEN_17237); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17832 = 6'h19 == state ? $signed(digest_39) : $signed(_GEN_17238); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17833 = 6'h19 == state ? $signed(digest_40) : $signed(_GEN_17239); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17834 = 6'h19 == state ? $signed(digest_41) : $signed(_GEN_17240); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17835 = 6'h19 == state ? $signed(digest_42) : $signed(_GEN_17241); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17836 = 6'h19 == state ? $signed(digest_43) : $signed(_GEN_17242); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17837 = 6'h19 == state ? $signed(digest_44) : $signed(_GEN_17243); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17838 = 6'h19 == state ? $signed(digest_45) : $signed(_GEN_17244); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17839 = 6'h19 == state ? $signed(digest_46) : $signed(_GEN_17245); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17840 = 6'h19 == state ? $signed(digest_47) : $signed(_GEN_17246); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17841 = 6'h19 == state ? $signed(digest_48) : $signed(_GEN_17247); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17842 = 6'h19 == state ? $signed(digest_49) : $signed(_GEN_17248); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17843 = 6'h19 == state ? $signed(digest_50) : $signed(_GEN_17249); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17844 = 6'h19 == state ? $signed(digest_51) : $signed(_GEN_17250); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17845 = 6'h19 == state ? $signed(digest_52) : $signed(_GEN_17251); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17846 = 6'h19 == state ? $signed(digest_53) : $signed(_GEN_17252); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17847 = 6'h19 == state ? $signed(digest_54) : $signed(_GEN_17253); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17848 = 6'h19 == state ? $signed(digest_55) : $signed(_GEN_17254); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17849 = 6'h19 == state ? $signed(digest_56) : $signed(_GEN_17255); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17850 = 6'h19 == state ? $signed(digest_57) : $signed(_GEN_17256); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17851 = 6'h19 == state ? $signed(digest_58) : $signed(_GEN_17257); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17852 = 6'h19 == state ? $signed(digest_59) : $signed(_GEN_17258); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17853 = 6'h19 == state ? $signed(digest_60) : $signed(_GEN_17259); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17854 = 6'h19 == state ? $signed(digest_61) : $signed(_GEN_17260); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17855 = 6'h19 == state ? $signed(digest_62) : $signed(_GEN_17261); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17856 = 6'h19 == state ? $signed(digest_63) : $signed(_GEN_17262); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17857 = 6'h19 == state ? $signed(digest_64) : $signed(_GEN_17263); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17858 = 6'h19 == state ? $signed(digest_65) : $signed(_GEN_17264); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17859 = 6'h19 == state ? $signed(digest_66) : $signed(_GEN_17265); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17860 = 6'h19 == state ? $signed(digest_67) : $signed(_GEN_17266); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17861 = 6'h19 == state ? $signed(digest_68) : $signed(_GEN_17267); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17862 = 6'h19 == state ? $signed(digest_69) : $signed(_GEN_17268); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17863 = 6'h19 == state ? $signed(digest_70) : $signed(_GEN_17269); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17864 = 6'h19 == state ? $signed(digest_71) : $signed(_GEN_17270); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17865 = 6'h19 == state ? $signed(digest_72) : $signed(_GEN_17271); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17866 = 6'h19 == state ? $signed(digest_73) : $signed(_GEN_17272); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17867 = 6'h19 == state ? $signed(digest_74) : $signed(_GEN_17273); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17868 = 6'h19 == state ? $signed(digest_75) : $signed(_GEN_17274); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17869 = 6'h19 == state ? $signed(digest_76) : $signed(_GEN_17275); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17870 = 6'h19 == state ? $signed(digest_77) : $signed(_GEN_17276); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17871 = 6'h19 == state ? $signed(digest_78) : $signed(_GEN_17277); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_17872 = 6'h19 == state ? $signed(digest_79) : $signed(_GEN_17278); // @[digest.scala 81:19 53:21]
  wire  _GEN_17874 = 6'h19 == state ? 1'h0 : _GEN_17280; // @[digest.scala 81:19 58:25]
  wire  _GEN_17957 = 6'h19 == state ? 1'h0 : _GEN_17363; // @[digest.scala 81:19 63:25]
  wire  _GEN_18040 = 6'h19 == state ? 1'h0 : _GEN_17446; // @[digest.scala 81:19 68:25]
  wire  _GEN_18123 = 6'h19 == state ? 1'h0 : _GEN_17529; // @[digest.scala 81:19 73:25]
  wire  _GEN_18206 = 6'h19 == state ? 1'h0 : _GEN_17612; // @[digest.scala 81:19 78:25]
  wire [5:0] _GEN_18207 = 6'h18 == state ? {{1'd0}, _state_T_8} : _GEN_17693; // @[digest.scala 179:19 81:19]
  wire [31:0] _GEN_18208 = 6'h18 == state ? $signed(w_0) : $signed(_GEN_17613); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18209 = 6'h18 == state ? $signed(w_1) : $signed(_GEN_17614); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18210 = 6'h18 == state ? $signed(w_2) : $signed(_GEN_17615); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18211 = 6'h18 == state ? $signed(w_3) : $signed(_GEN_17616); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18212 = 6'h18 == state ? $signed(w_4) : $signed(_GEN_17617); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18213 = 6'h18 == state ? $signed(w_5) : $signed(_GEN_17618); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18214 = 6'h18 == state ? $signed(w_6) : $signed(_GEN_17619); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18215 = 6'h18 == state ? $signed(w_7) : $signed(_GEN_17620); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18216 = 6'h18 == state ? $signed(w_8) : $signed(_GEN_17621); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18217 = 6'h18 == state ? $signed(w_9) : $signed(_GEN_17622); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18218 = 6'h18 == state ? $signed(w_10) : $signed(_GEN_17623); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18219 = 6'h18 == state ? $signed(w_11) : $signed(_GEN_17624); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18220 = 6'h18 == state ? $signed(w_12) : $signed(_GEN_17625); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18221 = 6'h18 == state ? $signed(w_13) : $signed(_GEN_17626); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18222 = 6'h18 == state ? $signed(w_14) : $signed(_GEN_17627); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18223 = 6'h18 == state ? $signed(w_15) : $signed(_GEN_17628); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18224 = 6'h18 == state ? $signed(w_16) : $signed(_GEN_17629); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18225 = 6'h18 == state ? $signed(w_17) : $signed(_GEN_17630); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18226 = 6'h18 == state ? $signed(w_18) : $signed(_GEN_17631); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18227 = 6'h18 == state ? $signed(w_19) : $signed(_GEN_17632); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18228 = 6'h18 == state ? $signed(w_20) : $signed(_GEN_17633); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18229 = 6'h18 == state ? $signed(w_21) : $signed(_GEN_17634); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18230 = 6'h18 == state ? $signed(w_22) : $signed(_GEN_17635); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18231 = 6'h18 == state ? $signed(w_23) : $signed(_GEN_17636); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18232 = 6'h18 == state ? $signed(w_24) : $signed(_GEN_17637); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18233 = 6'h18 == state ? $signed(w_25) : $signed(_GEN_17638); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18234 = 6'h18 == state ? $signed(w_26) : $signed(_GEN_17639); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18235 = 6'h18 == state ? $signed(w_27) : $signed(_GEN_17640); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18236 = 6'h18 == state ? $signed(w_28) : $signed(_GEN_17641); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18237 = 6'h18 == state ? $signed(w_29) : $signed(_GEN_17642); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18238 = 6'h18 == state ? $signed(w_30) : $signed(_GEN_17643); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18239 = 6'h18 == state ? $signed(w_31) : $signed(_GEN_17644); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18240 = 6'h18 == state ? $signed(w_32) : $signed(_GEN_17645); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18241 = 6'h18 == state ? $signed(w_33) : $signed(_GEN_17646); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18242 = 6'h18 == state ? $signed(w_34) : $signed(_GEN_17647); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18243 = 6'h18 == state ? $signed(w_35) : $signed(_GEN_17648); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18244 = 6'h18 == state ? $signed(w_36) : $signed(_GEN_17649); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18245 = 6'h18 == state ? $signed(w_37) : $signed(_GEN_17650); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18246 = 6'h18 == state ? $signed(w_38) : $signed(_GEN_17651); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18247 = 6'h18 == state ? $signed(w_39) : $signed(_GEN_17652); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18248 = 6'h18 == state ? $signed(w_40) : $signed(_GEN_17653); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18249 = 6'h18 == state ? $signed(w_41) : $signed(_GEN_17654); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18250 = 6'h18 == state ? $signed(w_42) : $signed(_GEN_17655); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18251 = 6'h18 == state ? $signed(w_43) : $signed(_GEN_17656); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18252 = 6'h18 == state ? $signed(w_44) : $signed(_GEN_17657); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18253 = 6'h18 == state ? $signed(w_45) : $signed(_GEN_17658); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18254 = 6'h18 == state ? $signed(w_46) : $signed(_GEN_17659); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18255 = 6'h18 == state ? $signed(w_47) : $signed(_GEN_17660); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18256 = 6'h18 == state ? $signed(w_48) : $signed(_GEN_17661); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18257 = 6'h18 == state ? $signed(w_49) : $signed(_GEN_17662); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18258 = 6'h18 == state ? $signed(w_50) : $signed(_GEN_17663); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18259 = 6'h18 == state ? $signed(w_51) : $signed(_GEN_17664); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18260 = 6'h18 == state ? $signed(w_52) : $signed(_GEN_17665); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18261 = 6'h18 == state ? $signed(w_53) : $signed(_GEN_17666); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18262 = 6'h18 == state ? $signed(w_54) : $signed(_GEN_17667); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18263 = 6'h18 == state ? $signed(w_55) : $signed(_GEN_17668); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18264 = 6'h18 == state ? $signed(w_56) : $signed(_GEN_17669); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18265 = 6'h18 == state ? $signed(w_57) : $signed(_GEN_17670); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18266 = 6'h18 == state ? $signed(w_58) : $signed(_GEN_17671); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18267 = 6'h18 == state ? $signed(w_59) : $signed(_GEN_17672); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18268 = 6'h18 == state ? $signed(w_60) : $signed(_GEN_17673); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18269 = 6'h18 == state ? $signed(w_61) : $signed(_GEN_17674); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18270 = 6'h18 == state ? $signed(w_62) : $signed(_GEN_17675); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18271 = 6'h18 == state ? $signed(w_63) : $signed(_GEN_17676); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18272 = 6'h18 == state ? $signed(w_64) : $signed(_GEN_17677); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18273 = 6'h18 == state ? $signed(w_65) : $signed(_GEN_17678); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18274 = 6'h18 == state ? $signed(w_66) : $signed(_GEN_17679); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18275 = 6'h18 == state ? $signed(w_67) : $signed(_GEN_17680); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18276 = 6'h18 == state ? $signed(w_68) : $signed(_GEN_17681); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18277 = 6'h18 == state ? $signed(w_69) : $signed(_GEN_17682); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18278 = 6'h18 == state ? $signed(w_70) : $signed(_GEN_17683); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18279 = 6'h18 == state ? $signed(w_71) : $signed(_GEN_17684); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18280 = 6'h18 == state ? $signed(w_72) : $signed(_GEN_17685); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18281 = 6'h18 == state ? $signed(w_73) : $signed(_GEN_17686); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18282 = 6'h18 == state ? $signed(w_74) : $signed(_GEN_17687); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18283 = 6'h18 == state ? $signed(w_75) : $signed(_GEN_17688); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18284 = 6'h18 == state ? $signed(w_76) : $signed(_GEN_17689); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18285 = 6'h18 == state ? $signed(w_77) : $signed(_GEN_17690); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18286 = 6'h18 == state ? $signed(w_78) : $signed(_GEN_17691); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18287 = 6'h18 == state ? $signed(w_79) : $signed(_GEN_17692); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18288 = 6'h18 == state ? $signed(temp) : $signed(_GEN_17694); // @[digest.scala 38:19 81:19]
  wire  _GEN_18289 = 6'h18 == state ? 1'h0 : _GEN_17695; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_18292 = 6'h18 == state ? $signed(t) : $signed(_GEN_17698); // @[digest.scala 35:16 81:19]
  wire  _GEN_18293 = 6'h18 == state ? 1'h0 : _GEN_17699; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_18296 = 6'h18 == state ? $signed(e) : $signed(_GEN_17702); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_18297 = 6'h18 == state ? $signed(d) : $signed(_GEN_17703); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_18298 = 6'h18 == state ? $signed(c) : $signed(_GEN_17704); // @[digest.scala 26:16 81:19]
  wire  _GEN_18299 = 6'h18 == state ? 1'h0 : _GEN_17705; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_18302 = 6'h18 == state ? $signed(b) : $signed(_GEN_17708); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_18303 = 6'h18 == state ? $signed(a) : $signed(_GEN_17709); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_18304 = 6'h18 == state ? $signed(j) : $signed(_GEN_17710); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_18305 = 6'h18 == state ? $signed(i) : $signed(_GEN_17711); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_18387 = 6'h18 == state ? $signed(digest_0) : $signed(_GEN_17793); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18388 = 6'h18 == state ? $signed(digest_1) : $signed(_GEN_17794); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18389 = 6'h18 == state ? $signed(digest_2) : $signed(_GEN_17795); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18390 = 6'h18 == state ? $signed(digest_3) : $signed(_GEN_17796); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18391 = 6'h18 == state ? $signed(digest_4) : $signed(_GEN_17797); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18392 = 6'h18 == state ? $signed(digest_5) : $signed(_GEN_17798); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18393 = 6'h18 == state ? $signed(digest_6) : $signed(_GEN_17799); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18394 = 6'h18 == state ? $signed(digest_7) : $signed(_GEN_17800); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18395 = 6'h18 == state ? $signed(digest_8) : $signed(_GEN_17801); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18396 = 6'h18 == state ? $signed(digest_9) : $signed(_GEN_17802); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18397 = 6'h18 == state ? $signed(digest_10) : $signed(_GEN_17803); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18398 = 6'h18 == state ? $signed(digest_11) : $signed(_GEN_17804); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18399 = 6'h18 == state ? $signed(digest_12) : $signed(_GEN_17805); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18400 = 6'h18 == state ? $signed(digest_13) : $signed(_GEN_17806); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18401 = 6'h18 == state ? $signed(digest_14) : $signed(_GEN_17807); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18402 = 6'h18 == state ? $signed(digest_15) : $signed(_GEN_17808); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18403 = 6'h18 == state ? $signed(digest_16) : $signed(_GEN_17809); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18404 = 6'h18 == state ? $signed(digest_17) : $signed(_GEN_17810); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18405 = 6'h18 == state ? $signed(digest_18) : $signed(_GEN_17811); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18406 = 6'h18 == state ? $signed(digest_19) : $signed(_GEN_17812); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18407 = 6'h18 == state ? $signed(digest_20) : $signed(_GEN_17813); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18408 = 6'h18 == state ? $signed(digest_21) : $signed(_GEN_17814); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18409 = 6'h18 == state ? $signed(digest_22) : $signed(_GEN_17815); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18410 = 6'h18 == state ? $signed(digest_23) : $signed(_GEN_17816); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18411 = 6'h18 == state ? $signed(digest_24) : $signed(_GEN_17817); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18412 = 6'h18 == state ? $signed(digest_25) : $signed(_GEN_17818); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18413 = 6'h18 == state ? $signed(digest_26) : $signed(_GEN_17819); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18414 = 6'h18 == state ? $signed(digest_27) : $signed(_GEN_17820); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18415 = 6'h18 == state ? $signed(digest_28) : $signed(_GEN_17821); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18416 = 6'h18 == state ? $signed(digest_29) : $signed(_GEN_17822); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18417 = 6'h18 == state ? $signed(digest_30) : $signed(_GEN_17823); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18418 = 6'h18 == state ? $signed(digest_31) : $signed(_GEN_17824); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18419 = 6'h18 == state ? $signed(digest_32) : $signed(_GEN_17825); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18420 = 6'h18 == state ? $signed(digest_33) : $signed(_GEN_17826); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18421 = 6'h18 == state ? $signed(digest_34) : $signed(_GEN_17827); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18422 = 6'h18 == state ? $signed(digest_35) : $signed(_GEN_17828); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18423 = 6'h18 == state ? $signed(digest_36) : $signed(_GEN_17829); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18424 = 6'h18 == state ? $signed(digest_37) : $signed(_GEN_17830); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18425 = 6'h18 == state ? $signed(digest_38) : $signed(_GEN_17831); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18426 = 6'h18 == state ? $signed(digest_39) : $signed(_GEN_17832); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18427 = 6'h18 == state ? $signed(digest_40) : $signed(_GEN_17833); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18428 = 6'h18 == state ? $signed(digest_41) : $signed(_GEN_17834); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18429 = 6'h18 == state ? $signed(digest_42) : $signed(_GEN_17835); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18430 = 6'h18 == state ? $signed(digest_43) : $signed(_GEN_17836); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18431 = 6'h18 == state ? $signed(digest_44) : $signed(_GEN_17837); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18432 = 6'h18 == state ? $signed(digest_45) : $signed(_GEN_17838); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18433 = 6'h18 == state ? $signed(digest_46) : $signed(_GEN_17839); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18434 = 6'h18 == state ? $signed(digest_47) : $signed(_GEN_17840); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18435 = 6'h18 == state ? $signed(digest_48) : $signed(_GEN_17841); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18436 = 6'h18 == state ? $signed(digest_49) : $signed(_GEN_17842); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18437 = 6'h18 == state ? $signed(digest_50) : $signed(_GEN_17843); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18438 = 6'h18 == state ? $signed(digest_51) : $signed(_GEN_17844); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18439 = 6'h18 == state ? $signed(digest_52) : $signed(_GEN_17845); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18440 = 6'h18 == state ? $signed(digest_53) : $signed(_GEN_17846); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18441 = 6'h18 == state ? $signed(digest_54) : $signed(_GEN_17847); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18442 = 6'h18 == state ? $signed(digest_55) : $signed(_GEN_17848); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18443 = 6'h18 == state ? $signed(digest_56) : $signed(_GEN_17849); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18444 = 6'h18 == state ? $signed(digest_57) : $signed(_GEN_17850); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18445 = 6'h18 == state ? $signed(digest_58) : $signed(_GEN_17851); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18446 = 6'h18 == state ? $signed(digest_59) : $signed(_GEN_17852); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18447 = 6'h18 == state ? $signed(digest_60) : $signed(_GEN_17853); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18448 = 6'h18 == state ? $signed(digest_61) : $signed(_GEN_17854); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18449 = 6'h18 == state ? $signed(digest_62) : $signed(_GEN_17855); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18450 = 6'h18 == state ? $signed(digest_63) : $signed(_GEN_17856); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18451 = 6'h18 == state ? $signed(digest_64) : $signed(_GEN_17857); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18452 = 6'h18 == state ? $signed(digest_65) : $signed(_GEN_17858); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18453 = 6'h18 == state ? $signed(digest_66) : $signed(_GEN_17859); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18454 = 6'h18 == state ? $signed(digest_67) : $signed(_GEN_17860); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18455 = 6'h18 == state ? $signed(digest_68) : $signed(_GEN_17861); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18456 = 6'h18 == state ? $signed(digest_69) : $signed(_GEN_17862); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18457 = 6'h18 == state ? $signed(digest_70) : $signed(_GEN_17863); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18458 = 6'h18 == state ? $signed(digest_71) : $signed(_GEN_17864); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18459 = 6'h18 == state ? $signed(digest_72) : $signed(_GEN_17865); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18460 = 6'h18 == state ? $signed(digest_73) : $signed(_GEN_17866); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18461 = 6'h18 == state ? $signed(digest_74) : $signed(_GEN_17867); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18462 = 6'h18 == state ? $signed(digest_75) : $signed(_GEN_17868); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18463 = 6'h18 == state ? $signed(digest_76) : $signed(_GEN_17869); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18464 = 6'h18 == state ? $signed(digest_77) : $signed(_GEN_17870); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18465 = 6'h18 == state ? $signed(digest_78) : $signed(_GEN_17871); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18466 = 6'h18 == state ? $signed(digest_79) : $signed(_GEN_17872); // @[digest.scala 81:19 53:21]
  wire  _GEN_18468 = 6'h18 == state ? 1'h0 : _GEN_17874; // @[digest.scala 81:19 58:25]
  wire  _GEN_18551 = 6'h18 == state ? 1'h0 : _GEN_17957; // @[digest.scala 81:19 63:25]
  wire  _GEN_18634 = 6'h18 == state ? 1'h0 : _GEN_18040; // @[digest.scala 81:19 68:25]
  wire  _GEN_18717 = 6'h18 == state ? 1'h0 : _GEN_18123; // @[digest.scala 81:19 73:25]
  wire  _GEN_18800 = 6'h18 == state ? 1'h0 : _GEN_18206; // @[digest.scala 81:19 78:25]
  wire [5:0] _GEN_18801 = 6'h17 == state ? _state_T_6 : _GEN_18207; // @[digest.scala 176:19 81:19]
  wire [31:0] _GEN_18802 = 6'h17 == state ? $signed(w_0) : $signed(_GEN_18208); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18803 = 6'h17 == state ? $signed(w_1) : $signed(_GEN_18209); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18804 = 6'h17 == state ? $signed(w_2) : $signed(_GEN_18210); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18805 = 6'h17 == state ? $signed(w_3) : $signed(_GEN_18211); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18806 = 6'h17 == state ? $signed(w_4) : $signed(_GEN_18212); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18807 = 6'h17 == state ? $signed(w_5) : $signed(_GEN_18213); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18808 = 6'h17 == state ? $signed(w_6) : $signed(_GEN_18214); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18809 = 6'h17 == state ? $signed(w_7) : $signed(_GEN_18215); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18810 = 6'h17 == state ? $signed(w_8) : $signed(_GEN_18216); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18811 = 6'h17 == state ? $signed(w_9) : $signed(_GEN_18217); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18812 = 6'h17 == state ? $signed(w_10) : $signed(_GEN_18218); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18813 = 6'h17 == state ? $signed(w_11) : $signed(_GEN_18219); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18814 = 6'h17 == state ? $signed(w_12) : $signed(_GEN_18220); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18815 = 6'h17 == state ? $signed(w_13) : $signed(_GEN_18221); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18816 = 6'h17 == state ? $signed(w_14) : $signed(_GEN_18222); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18817 = 6'h17 == state ? $signed(w_15) : $signed(_GEN_18223); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18818 = 6'h17 == state ? $signed(w_16) : $signed(_GEN_18224); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18819 = 6'h17 == state ? $signed(w_17) : $signed(_GEN_18225); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18820 = 6'h17 == state ? $signed(w_18) : $signed(_GEN_18226); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18821 = 6'h17 == state ? $signed(w_19) : $signed(_GEN_18227); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18822 = 6'h17 == state ? $signed(w_20) : $signed(_GEN_18228); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18823 = 6'h17 == state ? $signed(w_21) : $signed(_GEN_18229); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18824 = 6'h17 == state ? $signed(w_22) : $signed(_GEN_18230); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18825 = 6'h17 == state ? $signed(w_23) : $signed(_GEN_18231); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18826 = 6'h17 == state ? $signed(w_24) : $signed(_GEN_18232); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18827 = 6'h17 == state ? $signed(w_25) : $signed(_GEN_18233); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18828 = 6'h17 == state ? $signed(w_26) : $signed(_GEN_18234); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18829 = 6'h17 == state ? $signed(w_27) : $signed(_GEN_18235); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18830 = 6'h17 == state ? $signed(w_28) : $signed(_GEN_18236); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18831 = 6'h17 == state ? $signed(w_29) : $signed(_GEN_18237); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18832 = 6'h17 == state ? $signed(w_30) : $signed(_GEN_18238); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18833 = 6'h17 == state ? $signed(w_31) : $signed(_GEN_18239); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18834 = 6'h17 == state ? $signed(w_32) : $signed(_GEN_18240); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18835 = 6'h17 == state ? $signed(w_33) : $signed(_GEN_18241); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18836 = 6'h17 == state ? $signed(w_34) : $signed(_GEN_18242); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18837 = 6'h17 == state ? $signed(w_35) : $signed(_GEN_18243); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18838 = 6'h17 == state ? $signed(w_36) : $signed(_GEN_18244); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18839 = 6'h17 == state ? $signed(w_37) : $signed(_GEN_18245); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18840 = 6'h17 == state ? $signed(w_38) : $signed(_GEN_18246); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18841 = 6'h17 == state ? $signed(w_39) : $signed(_GEN_18247); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18842 = 6'h17 == state ? $signed(w_40) : $signed(_GEN_18248); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18843 = 6'h17 == state ? $signed(w_41) : $signed(_GEN_18249); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18844 = 6'h17 == state ? $signed(w_42) : $signed(_GEN_18250); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18845 = 6'h17 == state ? $signed(w_43) : $signed(_GEN_18251); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18846 = 6'h17 == state ? $signed(w_44) : $signed(_GEN_18252); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18847 = 6'h17 == state ? $signed(w_45) : $signed(_GEN_18253); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18848 = 6'h17 == state ? $signed(w_46) : $signed(_GEN_18254); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18849 = 6'h17 == state ? $signed(w_47) : $signed(_GEN_18255); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18850 = 6'h17 == state ? $signed(w_48) : $signed(_GEN_18256); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18851 = 6'h17 == state ? $signed(w_49) : $signed(_GEN_18257); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18852 = 6'h17 == state ? $signed(w_50) : $signed(_GEN_18258); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18853 = 6'h17 == state ? $signed(w_51) : $signed(_GEN_18259); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18854 = 6'h17 == state ? $signed(w_52) : $signed(_GEN_18260); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18855 = 6'h17 == state ? $signed(w_53) : $signed(_GEN_18261); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18856 = 6'h17 == state ? $signed(w_54) : $signed(_GEN_18262); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18857 = 6'h17 == state ? $signed(w_55) : $signed(_GEN_18263); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18858 = 6'h17 == state ? $signed(w_56) : $signed(_GEN_18264); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18859 = 6'h17 == state ? $signed(w_57) : $signed(_GEN_18265); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18860 = 6'h17 == state ? $signed(w_58) : $signed(_GEN_18266); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18861 = 6'h17 == state ? $signed(w_59) : $signed(_GEN_18267); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18862 = 6'h17 == state ? $signed(w_60) : $signed(_GEN_18268); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18863 = 6'h17 == state ? $signed(w_61) : $signed(_GEN_18269); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18864 = 6'h17 == state ? $signed(w_62) : $signed(_GEN_18270); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18865 = 6'h17 == state ? $signed(w_63) : $signed(_GEN_18271); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18866 = 6'h17 == state ? $signed(w_64) : $signed(_GEN_18272); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18867 = 6'h17 == state ? $signed(w_65) : $signed(_GEN_18273); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18868 = 6'h17 == state ? $signed(w_66) : $signed(_GEN_18274); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18869 = 6'h17 == state ? $signed(w_67) : $signed(_GEN_18275); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18870 = 6'h17 == state ? $signed(w_68) : $signed(_GEN_18276); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18871 = 6'h17 == state ? $signed(w_69) : $signed(_GEN_18277); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18872 = 6'h17 == state ? $signed(w_70) : $signed(_GEN_18278); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18873 = 6'h17 == state ? $signed(w_71) : $signed(_GEN_18279); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18874 = 6'h17 == state ? $signed(w_72) : $signed(_GEN_18280); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18875 = 6'h17 == state ? $signed(w_73) : $signed(_GEN_18281); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18876 = 6'h17 == state ? $signed(w_74) : $signed(_GEN_18282); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18877 = 6'h17 == state ? $signed(w_75) : $signed(_GEN_18283); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18878 = 6'h17 == state ? $signed(w_76) : $signed(_GEN_18284); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18879 = 6'h17 == state ? $signed(w_77) : $signed(_GEN_18285); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18880 = 6'h17 == state ? $signed(w_78) : $signed(_GEN_18286); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18881 = 6'h17 == state ? $signed(w_79) : $signed(_GEN_18287); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_18882 = 6'h17 == state ? $signed(temp) : $signed(_GEN_18288); // @[digest.scala 38:19 81:19]
  wire  _GEN_18883 = 6'h17 == state ? 1'h0 : _GEN_18289; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_18886 = 6'h17 == state ? $signed(t) : $signed(_GEN_18292); // @[digest.scala 35:16 81:19]
  wire  _GEN_18887 = 6'h17 == state ? 1'h0 : _GEN_18293; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_18890 = 6'h17 == state ? $signed(e) : $signed(_GEN_18296); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_18891 = 6'h17 == state ? $signed(d) : $signed(_GEN_18297); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_18892 = 6'h17 == state ? $signed(c) : $signed(_GEN_18298); // @[digest.scala 26:16 81:19]
  wire  _GEN_18893 = 6'h17 == state ? 1'h0 : _GEN_18299; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_18896 = 6'h17 == state ? $signed(b) : $signed(_GEN_18302); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_18897 = 6'h17 == state ? $signed(a) : $signed(_GEN_18303); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_18898 = 6'h17 == state ? $signed(j) : $signed(_GEN_18304); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_18899 = 6'h17 == state ? $signed(i) : $signed(_GEN_18305); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_18981 = 6'h17 == state ? $signed(digest_0) : $signed(_GEN_18387); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18982 = 6'h17 == state ? $signed(digest_1) : $signed(_GEN_18388); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18983 = 6'h17 == state ? $signed(digest_2) : $signed(_GEN_18389); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18984 = 6'h17 == state ? $signed(digest_3) : $signed(_GEN_18390); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18985 = 6'h17 == state ? $signed(digest_4) : $signed(_GEN_18391); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18986 = 6'h17 == state ? $signed(digest_5) : $signed(_GEN_18392); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18987 = 6'h17 == state ? $signed(digest_6) : $signed(_GEN_18393); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18988 = 6'h17 == state ? $signed(digest_7) : $signed(_GEN_18394); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18989 = 6'h17 == state ? $signed(digest_8) : $signed(_GEN_18395); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18990 = 6'h17 == state ? $signed(digest_9) : $signed(_GEN_18396); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18991 = 6'h17 == state ? $signed(digest_10) : $signed(_GEN_18397); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18992 = 6'h17 == state ? $signed(digest_11) : $signed(_GEN_18398); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18993 = 6'h17 == state ? $signed(digest_12) : $signed(_GEN_18399); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18994 = 6'h17 == state ? $signed(digest_13) : $signed(_GEN_18400); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18995 = 6'h17 == state ? $signed(digest_14) : $signed(_GEN_18401); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18996 = 6'h17 == state ? $signed(digest_15) : $signed(_GEN_18402); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18997 = 6'h17 == state ? $signed(digest_16) : $signed(_GEN_18403); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18998 = 6'h17 == state ? $signed(digest_17) : $signed(_GEN_18404); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_18999 = 6'h17 == state ? $signed(digest_18) : $signed(_GEN_18405); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19000 = 6'h17 == state ? $signed(digest_19) : $signed(_GEN_18406); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19001 = 6'h17 == state ? $signed(digest_20) : $signed(_GEN_18407); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19002 = 6'h17 == state ? $signed(digest_21) : $signed(_GEN_18408); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19003 = 6'h17 == state ? $signed(digest_22) : $signed(_GEN_18409); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19004 = 6'h17 == state ? $signed(digest_23) : $signed(_GEN_18410); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19005 = 6'h17 == state ? $signed(digest_24) : $signed(_GEN_18411); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19006 = 6'h17 == state ? $signed(digest_25) : $signed(_GEN_18412); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19007 = 6'h17 == state ? $signed(digest_26) : $signed(_GEN_18413); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19008 = 6'h17 == state ? $signed(digest_27) : $signed(_GEN_18414); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19009 = 6'h17 == state ? $signed(digest_28) : $signed(_GEN_18415); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19010 = 6'h17 == state ? $signed(digest_29) : $signed(_GEN_18416); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19011 = 6'h17 == state ? $signed(digest_30) : $signed(_GEN_18417); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19012 = 6'h17 == state ? $signed(digest_31) : $signed(_GEN_18418); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19013 = 6'h17 == state ? $signed(digest_32) : $signed(_GEN_18419); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19014 = 6'h17 == state ? $signed(digest_33) : $signed(_GEN_18420); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19015 = 6'h17 == state ? $signed(digest_34) : $signed(_GEN_18421); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19016 = 6'h17 == state ? $signed(digest_35) : $signed(_GEN_18422); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19017 = 6'h17 == state ? $signed(digest_36) : $signed(_GEN_18423); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19018 = 6'h17 == state ? $signed(digest_37) : $signed(_GEN_18424); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19019 = 6'h17 == state ? $signed(digest_38) : $signed(_GEN_18425); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19020 = 6'h17 == state ? $signed(digest_39) : $signed(_GEN_18426); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19021 = 6'h17 == state ? $signed(digest_40) : $signed(_GEN_18427); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19022 = 6'h17 == state ? $signed(digest_41) : $signed(_GEN_18428); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19023 = 6'h17 == state ? $signed(digest_42) : $signed(_GEN_18429); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19024 = 6'h17 == state ? $signed(digest_43) : $signed(_GEN_18430); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19025 = 6'h17 == state ? $signed(digest_44) : $signed(_GEN_18431); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19026 = 6'h17 == state ? $signed(digest_45) : $signed(_GEN_18432); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19027 = 6'h17 == state ? $signed(digest_46) : $signed(_GEN_18433); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19028 = 6'h17 == state ? $signed(digest_47) : $signed(_GEN_18434); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19029 = 6'h17 == state ? $signed(digest_48) : $signed(_GEN_18435); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19030 = 6'h17 == state ? $signed(digest_49) : $signed(_GEN_18436); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19031 = 6'h17 == state ? $signed(digest_50) : $signed(_GEN_18437); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19032 = 6'h17 == state ? $signed(digest_51) : $signed(_GEN_18438); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19033 = 6'h17 == state ? $signed(digest_52) : $signed(_GEN_18439); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19034 = 6'h17 == state ? $signed(digest_53) : $signed(_GEN_18440); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19035 = 6'h17 == state ? $signed(digest_54) : $signed(_GEN_18441); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19036 = 6'h17 == state ? $signed(digest_55) : $signed(_GEN_18442); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19037 = 6'h17 == state ? $signed(digest_56) : $signed(_GEN_18443); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19038 = 6'h17 == state ? $signed(digest_57) : $signed(_GEN_18444); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19039 = 6'h17 == state ? $signed(digest_58) : $signed(_GEN_18445); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19040 = 6'h17 == state ? $signed(digest_59) : $signed(_GEN_18446); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19041 = 6'h17 == state ? $signed(digest_60) : $signed(_GEN_18447); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19042 = 6'h17 == state ? $signed(digest_61) : $signed(_GEN_18448); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19043 = 6'h17 == state ? $signed(digest_62) : $signed(_GEN_18449); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19044 = 6'h17 == state ? $signed(digest_63) : $signed(_GEN_18450); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19045 = 6'h17 == state ? $signed(digest_64) : $signed(_GEN_18451); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19046 = 6'h17 == state ? $signed(digest_65) : $signed(_GEN_18452); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19047 = 6'h17 == state ? $signed(digest_66) : $signed(_GEN_18453); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19048 = 6'h17 == state ? $signed(digest_67) : $signed(_GEN_18454); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19049 = 6'h17 == state ? $signed(digest_68) : $signed(_GEN_18455); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19050 = 6'h17 == state ? $signed(digest_69) : $signed(_GEN_18456); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19051 = 6'h17 == state ? $signed(digest_70) : $signed(_GEN_18457); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19052 = 6'h17 == state ? $signed(digest_71) : $signed(_GEN_18458); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19053 = 6'h17 == state ? $signed(digest_72) : $signed(_GEN_18459); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19054 = 6'h17 == state ? $signed(digest_73) : $signed(_GEN_18460); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19055 = 6'h17 == state ? $signed(digest_74) : $signed(_GEN_18461); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19056 = 6'h17 == state ? $signed(digest_75) : $signed(_GEN_18462); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19057 = 6'h17 == state ? $signed(digest_76) : $signed(_GEN_18463); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19058 = 6'h17 == state ? $signed(digest_77) : $signed(_GEN_18464); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19059 = 6'h17 == state ? $signed(digest_78) : $signed(_GEN_18465); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19060 = 6'h17 == state ? $signed(digest_79) : $signed(_GEN_18466); // @[digest.scala 81:19 53:21]
  wire  _GEN_19062 = 6'h17 == state ? 1'h0 : _GEN_18468; // @[digest.scala 81:19 58:25]
  wire  _GEN_19145 = 6'h17 == state ? 1'h0 : _GEN_18551; // @[digest.scala 81:19 63:25]
  wire  _GEN_19228 = 6'h17 == state ? 1'h0 : _GEN_18634; // @[digest.scala 81:19 68:25]
  wire  _GEN_19311 = 6'h17 == state ? 1'h0 : _GEN_18717; // @[digest.scala 81:19 73:25]
  wire  _GEN_19394 = 6'h17 == state ? 1'h0 : _GEN_18800; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_19395 = 6'h16 == state ? $signed(32'sh0) : $signed(_GEN_18898); // @[digest.scala 172:15 81:19]
  wire [5:0] _GEN_19396 = 6'h16 == state ? 6'h17 : _GEN_18801; // @[digest.scala 173:19 81:19]
  wire [31:0] _GEN_19397 = 6'h16 == state ? $signed(w_0) : $signed(_GEN_18802); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19398 = 6'h16 == state ? $signed(w_1) : $signed(_GEN_18803); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19399 = 6'h16 == state ? $signed(w_2) : $signed(_GEN_18804); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19400 = 6'h16 == state ? $signed(w_3) : $signed(_GEN_18805); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19401 = 6'h16 == state ? $signed(w_4) : $signed(_GEN_18806); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19402 = 6'h16 == state ? $signed(w_5) : $signed(_GEN_18807); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19403 = 6'h16 == state ? $signed(w_6) : $signed(_GEN_18808); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19404 = 6'h16 == state ? $signed(w_7) : $signed(_GEN_18809); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19405 = 6'h16 == state ? $signed(w_8) : $signed(_GEN_18810); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19406 = 6'h16 == state ? $signed(w_9) : $signed(_GEN_18811); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19407 = 6'h16 == state ? $signed(w_10) : $signed(_GEN_18812); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19408 = 6'h16 == state ? $signed(w_11) : $signed(_GEN_18813); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19409 = 6'h16 == state ? $signed(w_12) : $signed(_GEN_18814); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19410 = 6'h16 == state ? $signed(w_13) : $signed(_GEN_18815); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19411 = 6'h16 == state ? $signed(w_14) : $signed(_GEN_18816); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19412 = 6'h16 == state ? $signed(w_15) : $signed(_GEN_18817); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19413 = 6'h16 == state ? $signed(w_16) : $signed(_GEN_18818); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19414 = 6'h16 == state ? $signed(w_17) : $signed(_GEN_18819); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19415 = 6'h16 == state ? $signed(w_18) : $signed(_GEN_18820); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19416 = 6'h16 == state ? $signed(w_19) : $signed(_GEN_18821); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19417 = 6'h16 == state ? $signed(w_20) : $signed(_GEN_18822); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19418 = 6'h16 == state ? $signed(w_21) : $signed(_GEN_18823); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19419 = 6'h16 == state ? $signed(w_22) : $signed(_GEN_18824); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19420 = 6'h16 == state ? $signed(w_23) : $signed(_GEN_18825); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19421 = 6'h16 == state ? $signed(w_24) : $signed(_GEN_18826); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19422 = 6'h16 == state ? $signed(w_25) : $signed(_GEN_18827); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19423 = 6'h16 == state ? $signed(w_26) : $signed(_GEN_18828); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19424 = 6'h16 == state ? $signed(w_27) : $signed(_GEN_18829); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19425 = 6'h16 == state ? $signed(w_28) : $signed(_GEN_18830); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19426 = 6'h16 == state ? $signed(w_29) : $signed(_GEN_18831); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19427 = 6'h16 == state ? $signed(w_30) : $signed(_GEN_18832); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19428 = 6'h16 == state ? $signed(w_31) : $signed(_GEN_18833); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19429 = 6'h16 == state ? $signed(w_32) : $signed(_GEN_18834); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19430 = 6'h16 == state ? $signed(w_33) : $signed(_GEN_18835); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19431 = 6'h16 == state ? $signed(w_34) : $signed(_GEN_18836); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19432 = 6'h16 == state ? $signed(w_35) : $signed(_GEN_18837); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19433 = 6'h16 == state ? $signed(w_36) : $signed(_GEN_18838); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19434 = 6'h16 == state ? $signed(w_37) : $signed(_GEN_18839); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19435 = 6'h16 == state ? $signed(w_38) : $signed(_GEN_18840); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19436 = 6'h16 == state ? $signed(w_39) : $signed(_GEN_18841); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19437 = 6'h16 == state ? $signed(w_40) : $signed(_GEN_18842); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19438 = 6'h16 == state ? $signed(w_41) : $signed(_GEN_18843); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19439 = 6'h16 == state ? $signed(w_42) : $signed(_GEN_18844); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19440 = 6'h16 == state ? $signed(w_43) : $signed(_GEN_18845); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19441 = 6'h16 == state ? $signed(w_44) : $signed(_GEN_18846); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19442 = 6'h16 == state ? $signed(w_45) : $signed(_GEN_18847); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19443 = 6'h16 == state ? $signed(w_46) : $signed(_GEN_18848); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19444 = 6'h16 == state ? $signed(w_47) : $signed(_GEN_18849); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19445 = 6'h16 == state ? $signed(w_48) : $signed(_GEN_18850); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19446 = 6'h16 == state ? $signed(w_49) : $signed(_GEN_18851); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19447 = 6'h16 == state ? $signed(w_50) : $signed(_GEN_18852); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19448 = 6'h16 == state ? $signed(w_51) : $signed(_GEN_18853); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19449 = 6'h16 == state ? $signed(w_52) : $signed(_GEN_18854); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19450 = 6'h16 == state ? $signed(w_53) : $signed(_GEN_18855); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19451 = 6'h16 == state ? $signed(w_54) : $signed(_GEN_18856); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19452 = 6'h16 == state ? $signed(w_55) : $signed(_GEN_18857); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19453 = 6'h16 == state ? $signed(w_56) : $signed(_GEN_18858); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19454 = 6'h16 == state ? $signed(w_57) : $signed(_GEN_18859); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19455 = 6'h16 == state ? $signed(w_58) : $signed(_GEN_18860); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19456 = 6'h16 == state ? $signed(w_59) : $signed(_GEN_18861); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19457 = 6'h16 == state ? $signed(w_60) : $signed(_GEN_18862); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19458 = 6'h16 == state ? $signed(w_61) : $signed(_GEN_18863); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19459 = 6'h16 == state ? $signed(w_62) : $signed(_GEN_18864); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19460 = 6'h16 == state ? $signed(w_63) : $signed(_GEN_18865); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19461 = 6'h16 == state ? $signed(w_64) : $signed(_GEN_18866); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19462 = 6'h16 == state ? $signed(w_65) : $signed(_GEN_18867); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19463 = 6'h16 == state ? $signed(w_66) : $signed(_GEN_18868); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19464 = 6'h16 == state ? $signed(w_67) : $signed(_GEN_18869); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19465 = 6'h16 == state ? $signed(w_68) : $signed(_GEN_18870); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19466 = 6'h16 == state ? $signed(w_69) : $signed(_GEN_18871); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19467 = 6'h16 == state ? $signed(w_70) : $signed(_GEN_18872); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19468 = 6'h16 == state ? $signed(w_71) : $signed(_GEN_18873); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19469 = 6'h16 == state ? $signed(w_72) : $signed(_GEN_18874); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19470 = 6'h16 == state ? $signed(w_73) : $signed(_GEN_18875); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19471 = 6'h16 == state ? $signed(w_74) : $signed(_GEN_18876); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19472 = 6'h16 == state ? $signed(w_75) : $signed(_GEN_18877); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19473 = 6'h16 == state ? $signed(w_76) : $signed(_GEN_18878); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19474 = 6'h16 == state ? $signed(w_77) : $signed(_GEN_18879); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19475 = 6'h16 == state ? $signed(w_78) : $signed(_GEN_18880); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19476 = 6'h16 == state ? $signed(w_79) : $signed(_GEN_18881); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19477 = 6'h16 == state ? $signed(temp) : $signed(_GEN_18882); // @[digest.scala 38:19 81:19]
  wire  _GEN_19478 = 6'h16 == state ? 1'h0 : _GEN_18883; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_19481 = 6'h16 == state ? $signed(t) : $signed(_GEN_18886); // @[digest.scala 35:16 81:19]
  wire  _GEN_19482 = 6'h16 == state ? 1'h0 : _GEN_18887; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_19485 = 6'h16 == state ? $signed(e) : $signed(_GEN_18890); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_19486 = 6'h16 == state ? $signed(d) : $signed(_GEN_18891); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_19487 = 6'h16 == state ? $signed(c) : $signed(_GEN_18892); // @[digest.scala 26:16 81:19]
  wire  _GEN_19488 = 6'h16 == state ? 1'h0 : _GEN_18893; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_19491 = 6'h16 == state ? $signed(b) : $signed(_GEN_18896); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_19492 = 6'h16 == state ? $signed(a) : $signed(_GEN_18897); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_19493 = 6'h16 == state ? $signed(i) : $signed(_GEN_18899); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_19575 = 6'h16 == state ? $signed(digest_0) : $signed(_GEN_18981); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19576 = 6'h16 == state ? $signed(digest_1) : $signed(_GEN_18982); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19577 = 6'h16 == state ? $signed(digest_2) : $signed(_GEN_18983); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19578 = 6'h16 == state ? $signed(digest_3) : $signed(_GEN_18984); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19579 = 6'h16 == state ? $signed(digest_4) : $signed(_GEN_18985); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19580 = 6'h16 == state ? $signed(digest_5) : $signed(_GEN_18986); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19581 = 6'h16 == state ? $signed(digest_6) : $signed(_GEN_18987); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19582 = 6'h16 == state ? $signed(digest_7) : $signed(_GEN_18988); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19583 = 6'h16 == state ? $signed(digest_8) : $signed(_GEN_18989); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19584 = 6'h16 == state ? $signed(digest_9) : $signed(_GEN_18990); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19585 = 6'h16 == state ? $signed(digest_10) : $signed(_GEN_18991); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19586 = 6'h16 == state ? $signed(digest_11) : $signed(_GEN_18992); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19587 = 6'h16 == state ? $signed(digest_12) : $signed(_GEN_18993); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19588 = 6'h16 == state ? $signed(digest_13) : $signed(_GEN_18994); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19589 = 6'h16 == state ? $signed(digest_14) : $signed(_GEN_18995); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19590 = 6'h16 == state ? $signed(digest_15) : $signed(_GEN_18996); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19591 = 6'h16 == state ? $signed(digest_16) : $signed(_GEN_18997); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19592 = 6'h16 == state ? $signed(digest_17) : $signed(_GEN_18998); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19593 = 6'h16 == state ? $signed(digest_18) : $signed(_GEN_18999); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19594 = 6'h16 == state ? $signed(digest_19) : $signed(_GEN_19000); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19595 = 6'h16 == state ? $signed(digest_20) : $signed(_GEN_19001); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19596 = 6'h16 == state ? $signed(digest_21) : $signed(_GEN_19002); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19597 = 6'h16 == state ? $signed(digest_22) : $signed(_GEN_19003); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19598 = 6'h16 == state ? $signed(digest_23) : $signed(_GEN_19004); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19599 = 6'h16 == state ? $signed(digest_24) : $signed(_GEN_19005); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19600 = 6'h16 == state ? $signed(digest_25) : $signed(_GEN_19006); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19601 = 6'h16 == state ? $signed(digest_26) : $signed(_GEN_19007); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19602 = 6'h16 == state ? $signed(digest_27) : $signed(_GEN_19008); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19603 = 6'h16 == state ? $signed(digest_28) : $signed(_GEN_19009); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19604 = 6'h16 == state ? $signed(digest_29) : $signed(_GEN_19010); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19605 = 6'h16 == state ? $signed(digest_30) : $signed(_GEN_19011); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19606 = 6'h16 == state ? $signed(digest_31) : $signed(_GEN_19012); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19607 = 6'h16 == state ? $signed(digest_32) : $signed(_GEN_19013); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19608 = 6'h16 == state ? $signed(digest_33) : $signed(_GEN_19014); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19609 = 6'h16 == state ? $signed(digest_34) : $signed(_GEN_19015); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19610 = 6'h16 == state ? $signed(digest_35) : $signed(_GEN_19016); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19611 = 6'h16 == state ? $signed(digest_36) : $signed(_GEN_19017); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19612 = 6'h16 == state ? $signed(digest_37) : $signed(_GEN_19018); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19613 = 6'h16 == state ? $signed(digest_38) : $signed(_GEN_19019); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19614 = 6'h16 == state ? $signed(digest_39) : $signed(_GEN_19020); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19615 = 6'h16 == state ? $signed(digest_40) : $signed(_GEN_19021); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19616 = 6'h16 == state ? $signed(digest_41) : $signed(_GEN_19022); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19617 = 6'h16 == state ? $signed(digest_42) : $signed(_GEN_19023); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19618 = 6'h16 == state ? $signed(digest_43) : $signed(_GEN_19024); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19619 = 6'h16 == state ? $signed(digest_44) : $signed(_GEN_19025); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19620 = 6'h16 == state ? $signed(digest_45) : $signed(_GEN_19026); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19621 = 6'h16 == state ? $signed(digest_46) : $signed(_GEN_19027); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19622 = 6'h16 == state ? $signed(digest_47) : $signed(_GEN_19028); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19623 = 6'h16 == state ? $signed(digest_48) : $signed(_GEN_19029); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19624 = 6'h16 == state ? $signed(digest_49) : $signed(_GEN_19030); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19625 = 6'h16 == state ? $signed(digest_50) : $signed(_GEN_19031); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19626 = 6'h16 == state ? $signed(digest_51) : $signed(_GEN_19032); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19627 = 6'h16 == state ? $signed(digest_52) : $signed(_GEN_19033); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19628 = 6'h16 == state ? $signed(digest_53) : $signed(_GEN_19034); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19629 = 6'h16 == state ? $signed(digest_54) : $signed(_GEN_19035); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19630 = 6'h16 == state ? $signed(digest_55) : $signed(_GEN_19036); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19631 = 6'h16 == state ? $signed(digest_56) : $signed(_GEN_19037); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19632 = 6'h16 == state ? $signed(digest_57) : $signed(_GEN_19038); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19633 = 6'h16 == state ? $signed(digest_58) : $signed(_GEN_19039); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19634 = 6'h16 == state ? $signed(digest_59) : $signed(_GEN_19040); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19635 = 6'h16 == state ? $signed(digest_60) : $signed(_GEN_19041); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19636 = 6'h16 == state ? $signed(digest_61) : $signed(_GEN_19042); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19637 = 6'h16 == state ? $signed(digest_62) : $signed(_GEN_19043); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19638 = 6'h16 == state ? $signed(digest_63) : $signed(_GEN_19044); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19639 = 6'h16 == state ? $signed(digest_64) : $signed(_GEN_19045); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19640 = 6'h16 == state ? $signed(digest_65) : $signed(_GEN_19046); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19641 = 6'h16 == state ? $signed(digest_66) : $signed(_GEN_19047); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19642 = 6'h16 == state ? $signed(digest_67) : $signed(_GEN_19048); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19643 = 6'h16 == state ? $signed(digest_68) : $signed(_GEN_19049); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19644 = 6'h16 == state ? $signed(digest_69) : $signed(_GEN_19050); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19645 = 6'h16 == state ? $signed(digest_70) : $signed(_GEN_19051); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19646 = 6'h16 == state ? $signed(digest_71) : $signed(_GEN_19052); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19647 = 6'h16 == state ? $signed(digest_72) : $signed(_GEN_19053); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19648 = 6'h16 == state ? $signed(digest_73) : $signed(_GEN_19054); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19649 = 6'h16 == state ? $signed(digest_74) : $signed(_GEN_19055); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19650 = 6'h16 == state ? $signed(digest_75) : $signed(_GEN_19056); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19651 = 6'h16 == state ? $signed(digest_76) : $signed(_GEN_19057); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19652 = 6'h16 == state ? $signed(digest_77) : $signed(_GEN_19058); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19653 = 6'h16 == state ? $signed(digest_78) : $signed(_GEN_19059); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_19654 = 6'h16 == state ? $signed(digest_79) : $signed(_GEN_19060); // @[digest.scala 81:19 53:21]
  wire  _GEN_19656 = 6'h16 == state ? 1'h0 : _GEN_19062; // @[digest.scala 81:19 58:25]
  wire  _GEN_19739 = 6'h16 == state ? 1'h0 : _GEN_19145; // @[digest.scala 81:19 63:25]
  wire  _GEN_19822 = 6'h16 == state ? 1'h0 : _GEN_19228; // @[digest.scala 81:19 68:25]
  wire  _GEN_19905 = 6'h16 == state ? 1'h0 : _GEN_19311; // @[digest.scala 81:19 73:25]
  wire  _GEN_19988 = 6'h16 == state ? 1'h0 : _GEN_19394; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_19989 = 6'h15 == state ? $signed(e) : $signed(olde); // @[digest.scala 168:18 33:19 81:19]
  wire [5:0] _GEN_19990 = 6'h15 == state ? 6'h16 : _GEN_19396; // @[digest.scala 169:19 81:19]
  wire [31:0] _GEN_19991 = 6'h15 == state ? $signed(j) : $signed(_GEN_19395); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_19992 = 6'h15 == state ? $signed(w_0) : $signed(_GEN_19397); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19993 = 6'h15 == state ? $signed(w_1) : $signed(_GEN_19398); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19994 = 6'h15 == state ? $signed(w_2) : $signed(_GEN_19399); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19995 = 6'h15 == state ? $signed(w_3) : $signed(_GEN_19400); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19996 = 6'h15 == state ? $signed(w_4) : $signed(_GEN_19401); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19997 = 6'h15 == state ? $signed(w_5) : $signed(_GEN_19402); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19998 = 6'h15 == state ? $signed(w_6) : $signed(_GEN_19403); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_19999 = 6'h15 == state ? $signed(w_7) : $signed(_GEN_19404); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20000 = 6'h15 == state ? $signed(w_8) : $signed(_GEN_19405); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20001 = 6'h15 == state ? $signed(w_9) : $signed(_GEN_19406); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20002 = 6'h15 == state ? $signed(w_10) : $signed(_GEN_19407); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20003 = 6'h15 == state ? $signed(w_11) : $signed(_GEN_19408); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20004 = 6'h15 == state ? $signed(w_12) : $signed(_GEN_19409); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20005 = 6'h15 == state ? $signed(w_13) : $signed(_GEN_19410); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20006 = 6'h15 == state ? $signed(w_14) : $signed(_GEN_19411); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20007 = 6'h15 == state ? $signed(w_15) : $signed(_GEN_19412); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20008 = 6'h15 == state ? $signed(w_16) : $signed(_GEN_19413); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20009 = 6'h15 == state ? $signed(w_17) : $signed(_GEN_19414); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20010 = 6'h15 == state ? $signed(w_18) : $signed(_GEN_19415); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20011 = 6'h15 == state ? $signed(w_19) : $signed(_GEN_19416); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20012 = 6'h15 == state ? $signed(w_20) : $signed(_GEN_19417); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20013 = 6'h15 == state ? $signed(w_21) : $signed(_GEN_19418); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20014 = 6'h15 == state ? $signed(w_22) : $signed(_GEN_19419); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20015 = 6'h15 == state ? $signed(w_23) : $signed(_GEN_19420); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20016 = 6'h15 == state ? $signed(w_24) : $signed(_GEN_19421); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20017 = 6'h15 == state ? $signed(w_25) : $signed(_GEN_19422); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20018 = 6'h15 == state ? $signed(w_26) : $signed(_GEN_19423); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20019 = 6'h15 == state ? $signed(w_27) : $signed(_GEN_19424); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20020 = 6'h15 == state ? $signed(w_28) : $signed(_GEN_19425); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20021 = 6'h15 == state ? $signed(w_29) : $signed(_GEN_19426); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20022 = 6'h15 == state ? $signed(w_30) : $signed(_GEN_19427); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20023 = 6'h15 == state ? $signed(w_31) : $signed(_GEN_19428); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20024 = 6'h15 == state ? $signed(w_32) : $signed(_GEN_19429); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20025 = 6'h15 == state ? $signed(w_33) : $signed(_GEN_19430); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20026 = 6'h15 == state ? $signed(w_34) : $signed(_GEN_19431); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20027 = 6'h15 == state ? $signed(w_35) : $signed(_GEN_19432); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20028 = 6'h15 == state ? $signed(w_36) : $signed(_GEN_19433); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20029 = 6'h15 == state ? $signed(w_37) : $signed(_GEN_19434); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20030 = 6'h15 == state ? $signed(w_38) : $signed(_GEN_19435); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20031 = 6'h15 == state ? $signed(w_39) : $signed(_GEN_19436); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20032 = 6'h15 == state ? $signed(w_40) : $signed(_GEN_19437); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20033 = 6'h15 == state ? $signed(w_41) : $signed(_GEN_19438); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20034 = 6'h15 == state ? $signed(w_42) : $signed(_GEN_19439); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20035 = 6'h15 == state ? $signed(w_43) : $signed(_GEN_19440); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20036 = 6'h15 == state ? $signed(w_44) : $signed(_GEN_19441); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20037 = 6'h15 == state ? $signed(w_45) : $signed(_GEN_19442); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20038 = 6'h15 == state ? $signed(w_46) : $signed(_GEN_19443); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20039 = 6'h15 == state ? $signed(w_47) : $signed(_GEN_19444); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20040 = 6'h15 == state ? $signed(w_48) : $signed(_GEN_19445); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20041 = 6'h15 == state ? $signed(w_49) : $signed(_GEN_19446); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20042 = 6'h15 == state ? $signed(w_50) : $signed(_GEN_19447); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20043 = 6'h15 == state ? $signed(w_51) : $signed(_GEN_19448); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20044 = 6'h15 == state ? $signed(w_52) : $signed(_GEN_19449); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20045 = 6'h15 == state ? $signed(w_53) : $signed(_GEN_19450); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20046 = 6'h15 == state ? $signed(w_54) : $signed(_GEN_19451); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20047 = 6'h15 == state ? $signed(w_55) : $signed(_GEN_19452); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20048 = 6'h15 == state ? $signed(w_56) : $signed(_GEN_19453); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20049 = 6'h15 == state ? $signed(w_57) : $signed(_GEN_19454); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20050 = 6'h15 == state ? $signed(w_58) : $signed(_GEN_19455); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20051 = 6'h15 == state ? $signed(w_59) : $signed(_GEN_19456); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20052 = 6'h15 == state ? $signed(w_60) : $signed(_GEN_19457); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20053 = 6'h15 == state ? $signed(w_61) : $signed(_GEN_19458); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20054 = 6'h15 == state ? $signed(w_62) : $signed(_GEN_19459); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20055 = 6'h15 == state ? $signed(w_63) : $signed(_GEN_19460); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20056 = 6'h15 == state ? $signed(w_64) : $signed(_GEN_19461); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20057 = 6'h15 == state ? $signed(w_65) : $signed(_GEN_19462); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20058 = 6'h15 == state ? $signed(w_66) : $signed(_GEN_19463); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20059 = 6'h15 == state ? $signed(w_67) : $signed(_GEN_19464); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20060 = 6'h15 == state ? $signed(w_68) : $signed(_GEN_19465); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20061 = 6'h15 == state ? $signed(w_69) : $signed(_GEN_19466); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20062 = 6'h15 == state ? $signed(w_70) : $signed(_GEN_19467); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20063 = 6'h15 == state ? $signed(w_71) : $signed(_GEN_19468); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20064 = 6'h15 == state ? $signed(w_72) : $signed(_GEN_19469); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20065 = 6'h15 == state ? $signed(w_73) : $signed(_GEN_19470); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20066 = 6'h15 == state ? $signed(w_74) : $signed(_GEN_19471); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20067 = 6'h15 == state ? $signed(w_75) : $signed(_GEN_19472); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20068 = 6'h15 == state ? $signed(w_76) : $signed(_GEN_19473); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20069 = 6'h15 == state ? $signed(w_77) : $signed(_GEN_19474); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20070 = 6'h15 == state ? $signed(w_78) : $signed(_GEN_19475); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20071 = 6'h15 == state ? $signed(w_79) : $signed(_GEN_19476); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20072 = 6'h15 == state ? $signed(temp) : $signed(_GEN_19477); // @[digest.scala 38:19 81:19]
  wire  _GEN_20073 = 6'h15 == state ? 1'h0 : _GEN_19478; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_20076 = 6'h15 == state ? $signed(t) : $signed(_GEN_19481); // @[digest.scala 35:16 81:19]
  wire  _GEN_20077 = 6'h15 == state ? 1'h0 : _GEN_19482; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_20080 = 6'h15 == state ? $signed(e) : $signed(_GEN_19485); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_20081 = 6'h15 == state ? $signed(d) : $signed(_GEN_19486); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_20082 = 6'h15 == state ? $signed(c) : $signed(_GEN_19487); // @[digest.scala 26:16 81:19]
  wire  _GEN_20083 = 6'h15 == state ? 1'h0 : _GEN_19488; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_20086 = 6'h15 == state ? $signed(b) : $signed(_GEN_19491); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_20087 = 6'h15 == state ? $signed(a) : $signed(_GEN_19492); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_20088 = 6'h15 == state ? $signed(i) : $signed(_GEN_19493); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_20170 = 6'h15 == state ? $signed(digest_0) : $signed(_GEN_19575); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20171 = 6'h15 == state ? $signed(digest_1) : $signed(_GEN_19576); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20172 = 6'h15 == state ? $signed(digest_2) : $signed(_GEN_19577); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20173 = 6'h15 == state ? $signed(digest_3) : $signed(_GEN_19578); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20174 = 6'h15 == state ? $signed(digest_4) : $signed(_GEN_19579); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20175 = 6'h15 == state ? $signed(digest_5) : $signed(_GEN_19580); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20176 = 6'h15 == state ? $signed(digest_6) : $signed(_GEN_19581); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20177 = 6'h15 == state ? $signed(digest_7) : $signed(_GEN_19582); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20178 = 6'h15 == state ? $signed(digest_8) : $signed(_GEN_19583); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20179 = 6'h15 == state ? $signed(digest_9) : $signed(_GEN_19584); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20180 = 6'h15 == state ? $signed(digest_10) : $signed(_GEN_19585); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20181 = 6'h15 == state ? $signed(digest_11) : $signed(_GEN_19586); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20182 = 6'h15 == state ? $signed(digest_12) : $signed(_GEN_19587); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20183 = 6'h15 == state ? $signed(digest_13) : $signed(_GEN_19588); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20184 = 6'h15 == state ? $signed(digest_14) : $signed(_GEN_19589); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20185 = 6'h15 == state ? $signed(digest_15) : $signed(_GEN_19590); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20186 = 6'h15 == state ? $signed(digest_16) : $signed(_GEN_19591); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20187 = 6'h15 == state ? $signed(digest_17) : $signed(_GEN_19592); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20188 = 6'h15 == state ? $signed(digest_18) : $signed(_GEN_19593); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20189 = 6'h15 == state ? $signed(digest_19) : $signed(_GEN_19594); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20190 = 6'h15 == state ? $signed(digest_20) : $signed(_GEN_19595); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20191 = 6'h15 == state ? $signed(digest_21) : $signed(_GEN_19596); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20192 = 6'h15 == state ? $signed(digest_22) : $signed(_GEN_19597); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20193 = 6'h15 == state ? $signed(digest_23) : $signed(_GEN_19598); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20194 = 6'h15 == state ? $signed(digest_24) : $signed(_GEN_19599); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20195 = 6'h15 == state ? $signed(digest_25) : $signed(_GEN_19600); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20196 = 6'h15 == state ? $signed(digest_26) : $signed(_GEN_19601); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20197 = 6'h15 == state ? $signed(digest_27) : $signed(_GEN_19602); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20198 = 6'h15 == state ? $signed(digest_28) : $signed(_GEN_19603); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20199 = 6'h15 == state ? $signed(digest_29) : $signed(_GEN_19604); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20200 = 6'h15 == state ? $signed(digest_30) : $signed(_GEN_19605); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20201 = 6'h15 == state ? $signed(digest_31) : $signed(_GEN_19606); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20202 = 6'h15 == state ? $signed(digest_32) : $signed(_GEN_19607); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20203 = 6'h15 == state ? $signed(digest_33) : $signed(_GEN_19608); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20204 = 6'h15 == state ? $signed(digest_34) : $signed(_GEN_19609); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20205 = 6'h15 == state ? $signed(digest_35) : $signed(_GEN_19610); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20206 = 6'h15 == state ? $signed(digest_36) : $signed(_GEN_19611); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20207 = 6'h15 == state ? $signed(digest_37) : $signed(_GEN_19612); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20208 = 6'h15 == state ? $signed(digest_38) : $signed(_GEN_19613); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20209 = 6'h15 == state ? $signed(digest_39) : $signed(_GEN_19614); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20210 = 6'h15 == state ? $signed(digest_40) : $signed(_GEN_19615); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20211 = 6'h15 == state ? $signed(digest_41) : $signed(_GEN_19616); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20212 = 6'h15 == state ? $signed(digest_42) : $signed(_GEN_19617); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20213 = 6'h15 == state ? $signed(digest_43) : $signed(_GEN_19618); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20214 = 6'h15 == state ? $signed(digest_44) : $signed(_GEN_19619); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20215 = 6'h15 == state ? $signed(digest_45) : $signed(_GEN_19620); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20216 = 6'h15 == state ? $signed(digest_46) : $signed(_GEN_19621); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20217 = 6'h15 == state ? $signed(digest_47) : $signed(_GEN_19622); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20218 = 6'h15 == state ? $signed(digest_48) : $signed(_GEN_19623); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20219 = 6'h15 == state ? $signed(digest_49) : $signed(_GEN_19624); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20220 = 6'h15 == state ? $signed(digest_50) : $signed(_GEN_19625); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20221 = 6'h15 == state ? $signed(digest_51) : $signed(_GEN_19626); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20222 = 6'h15 == state ? $signed(digest_52) : $signed(_GEN_19627); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20223 = 6'h15 == state ? $signed(digest_53) : $signed(_GEN_19628); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20224 = 6'h15 == state ? $signed(digest_54) : $signed(_GEN_19629); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20225 = 6'h15 == state ? $signed(digest_55) : $signed(_GEN_19630); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20226 = 6'h15 == state ? $signed(digest_56) : $signed(_GEN_19631); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20227 = 6'h15 == state ? $signed(digest_57) : $signed(_GEN_19632); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20228 = 6'h15 == state ? $signed(digest_58) : $signed(_GEN_19633); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20229 = 6'h15 == state ? $signed(digest_59) : $signed(_GEN_19634); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20230 = 6'h15 == state ? $signed(digest_60) : $signed(_GEN_19635); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20231 = 6'h15 == state ? $signed(digest_61) : $signed(_GEN_19636); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20232 = 6'h15 == state ? $signed(digest_62) : $signed(_GEN_19637); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20233 = 6'h15 == state ? $signed(digest_63) : $signed(_GEN_19638); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20234 = 6'h15 == state ? $signed(digest_64) : $signed(_GEN_19639); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20235 = 6'h15 == state ? $signed(digest_65) : $signed(_GEN_19640); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20236 = 6'h15 == state ? $signed(digest_66) : $signed(_GEN_19641); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20237 = 6'h15 == state ? $signed(digest_67) : $signed(_GEN_19642); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20238 = 6'h15 == state ? $signed(digest_68) : $signed(_GEN_19643); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20239 = 6'h15 == state ? $signed(digest_69) : $signed(_GEN_19644); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20240 = 6'h15 == state ? $signed(digest_70) : $signed(_GEN_19645); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20241 = 6'h15 == state ? $signed(digest_71) : $signed(_GEN_19646); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20242 = 6'h15 == state ? $signed(digest_72) : $signed(_GEN_19647); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20243 = 6'h15 == state ? $signed(digest_73) : $signed(_GEN_19648); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20244 = 6'h15 == state ? $signed(digest_74) : $signed(_GEN_19649); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20245 = 6'h15 == state ? $signed(digest_75) : $signed(_GEN_19650); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20246 = 6'h15 == state ? $signed(digest_76) : $signed(_GEN_19651); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20247 = 6'h15 == state ? $signed(digest_77) : $signed(_GEN_19652); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20248 = 6'h15 == state ? $signed(digest_78) : $signed(_GEN_19653); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20249 = 6'h15 == state ? $signed(digest_79) : $signed(_GEN_19654); // @[digest.scala 81:19 53:21]
  wire  _GEN_20251 = 6'h15 == state ? 1'h0 : _GEN_19656; // @[digest.scala 81:19 58:25]
  wire  _GEN_20334 = 6'h15 == state ? 1'h0 : _GEN_19739; // @[digest.scala 81:19 63:25]
  wire  _GEN_20417 = 6'h15 == state ? 1'h0 : _GEN_19822; // @[digest.scala 81:19 68:25]
  wire  _GEN_20500 = 6'h15 == state ? 1'h0 : _GEN_19905; // @[digest.scala 81:19 73:25]
  wire  _GEN_20583 = 6'h15 == state ? 1'h0 : _GEN_19988; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_20584 = 6'h14 == state ? $signed(d) : $signed(oldd); // @[digest.scala 164:18 32:19 81:19]
  wire [5:0] _GEN_20585 = 6'h14 == state ? 6'h15 : _GEN_19990; // @[digest.scala 165:19 81:19]
  wire [31:0] _GEN_20586 = 6'h14 == state ? $signed(olde) : $signed(_GEN_19989); // @[digest.scala 33:19 81:19]
  wire [31:0] _GEN_20587 = 6'h14 == state ? $signed(j) : $signed(_GEN_19991); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_20588 = 6'h14 == state ? $signed(w_0) : $signed(_GEN_19992); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20589 = 6'h14 == state ? $signed(w_1) : $signed(_GEN_19993); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20590 = 6'h14 == state ? $signed(w_2) : $signed(_GEN_19994); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20591 = 6'h14 == state ? $signed(w_3) : $signed(_GEN_19995); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20592 = 6'h14 == state ? $signed(w_4) : $signed(_GEN_19996); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20593 = 6'h14 == state ? $signed(w_5) : $signed(_GEN_19997); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20594 = 6'h14 == state ? $signed(w_6) : $signed(_GEN_19998); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20595 = 6'h14 == state ? $signed(w_7) : $signed(_GEN_19999); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20596 = 6'h14 == state ? $signed(w_8) : $signed(_GEN_20000); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20597 = 6'h14 == state ? $signed(w_9) : $signed(_GEN_20001); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20598 = 6'h14 == state ? $signed(w_10) : $signed(_GEN_20002); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20599 = 6'h14 == state ? $signed(w_11) : $signed(_GEN_20003); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20600 = 6'h14 == state ? $signed(w_12) : $signed(_GEN_20004); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20601 = 6'h14 == state ? $signed(w_13) : $signed(_GEN_20005); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20602 = 6'h14 == state ? $signed(w_14) : $signed(_GEN_20006); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20603 = 6'h14 == state ? $signed(w_15) : $signed(_GEN_20007); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20604 = 6'h14 == state ? $signed(w_16) : $signed(_GEN_20008); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20605 = 6'h14 == state ? $signed(w_17) : $signed(_GEN_20009); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20606 = 6'h14 == state ? $signed(w_18) : $signed(_GEN_20010); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20607 = 6'h14 == state ? $signed(w_19) : $signed(_GEN_20011); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20608 = 6'h14 == state ? $signed(w_20) : $signed(_GEN_20012); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20609 = 6'h14 == state ? $signed(w_21) : $signed(_GEN_20013); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20610 = 6'h14 == state ? $signed(w_22) : $signed(_GEN_20014); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20611 = 6'h14 == state ? $signed(w_23) : $signed(_GEN_20015); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20612 = 6'h14 == state ? $signed(w_24) : $signed(_GEN_20016); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20613 = 6'h14 == state ? $signed(w_25) : $signed(_GEN_20017); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20614 = 6'h14 == state ? $signed(w_26) : $signed(_GEN_20018); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20615 = 6'h14 == state ? $signed(w_27) : $signed(_GEN_20019); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20616 = 6'h14 == state ? $signed(w_28) : $signed(_GEN_20020); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20617 = 6'h14 == state ? $signed(w_29) : $signed(_GEN_20021); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20618 = 6'h14 == state ? $signed(w_30) : $signed(_GEN_20022); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20619 = 6'h14 == state ? $signed(w_31) : $signed(_GEN_20023); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20620 = 6'h14 == state ? $signed(w_32) : $signed(_GEN_20024); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20621 = 6'h14 == state ? $signed(w_33) : $signed(_GEN_20025); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20622 = 6'h14 == state ? $signed(w_34) : $signed(_GEN_20026); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20623 = 6'h14 == state ? $signed(w_35) : $signed(_GEN_20027); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20624 = 6'h14 == state ? $signed(w_36) : $signed(_GEN_20028); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20625 = 6'h14 == state ? $signed(w_37) : $signed(_GEN_20029); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20626 = 6'h14 == state ? $signed(w_38) : $signed(_GEN_20030); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20627 = 6'h14 == state ? $signed(w_39) : $signed(_GEN_20031); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20628 = 6'h14 == state ? $signed(w_40) : $signed(_GEN_20032); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20629 = 6'h14 == state ? $signed(w_41) : $signed(_GEN_20033); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20630 = 6'h14 == state ? $signed(w_42) : $signed(_GEN_20034); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20631 = 6'h14 == state ? $signed(w_43) : $signed(_GEN_20035); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20632 = 6'h14 == state ? $signed(w_44) : $signed(_GEN_20036); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20633 = 6'h14 == state ? $signed(w_45) : $signed(_GEN_20037); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20634 = 6'h14 == state ? $signed(w_46) : $signed(_GEN_20038); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20635 = 6'h14 == state ? $signed(w_47) : $signed(_GEN_20039); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20636 = 6'h14 == state ? $signed(w_48) : $signed(_GEN_20040); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20637 = 6'h14 == state ? $signed(w_49) : $signed(_GEN_20041); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20638 = 6'h14 == state ? $signed(w_50) : $signed(_GEN_20042); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20639 = 6'h14 == state ? $signed(w_51) : $signed(_GEN_20043); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20640 = 6'h14 == state ? $signed(w_52) : $signed(_GEN_20044); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20641 = 6'h14 == state ? $signed(w_53) : $signed(_GEN_20045); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20642 = 6'h14 == state ? $signed(w_54) : $signed(_GEN_20046); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20643 = 6'h14 == state ? $signed(w_55) : $signed(_GEN_20047); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20644 = 6'h14 == state ? $signed(w_56) : $signed(_GEN_20048); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20645 = 6'h14 == state ? $signed(w_57) : $signed(_GEN_20049); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20646 = 6'h14 == state ? $signed(w_58) : $signed(_GEN_20050); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20647 = 6'h14 == state ? $signed(w_59) : $signed(_GEN_20051); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20648 = 6'h14 == state ? $signed(w_60) : $signed(_GEN_20052); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20649 = 6'h14 == state ? $signed(w_61) : $signed(_GEN_20053); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20650 = 6'h14 == state ? $signed(w_62) : $signed(_GEN_20054); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20651 = 6'h14 == state ? $signed(w_63) : $signed(_GEN_20055); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20652 = 6'h14 == state ? $signed(w_64) : $signed(_GEN_20056); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20653 = 6'h14 == state ? $signed(w_65) : $signed(_GEN_20057); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20654 = 6'h14 == state ? $signed(w_66) : $signed(_GEN_20058); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20655 = 6'h14 == state ? $signed(w_67) : $signed(_GEN_20059); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20656 = 6'h14 == state ? $signed(w_68) : $signed(_GEN_20060); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20657 = 6'h14 == state ? $signed(w_69) : $signed(_GEN_20061); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20658 = 6'h14 == state ? $signed(w_70) : $signed(_GEN_20062); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20659 = 6'h14 == state ? $signed(w_71) : $signed(_GEN_20063); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20660 = 6'h14 == state ? $signed(w_72) : $signed(_GEN_20064); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20661 = 6'h14 == state ? $signed(w_73) : $signed(_GEN_20065); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20662 = 6'h14 == state ? $signed(w_74) : $signed(_GEN_20066); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20663 = 6'h14 == state ? $signed(w_75) : $signed(_GEN_20067); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20664 = 6'h14 == state ? $signed(w_76) : $signed(_GEN_20068); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20665 = 6'h14 == state ? $signed(w_77) : $signed(_GEN_20069); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20666 = 6'h14 == state ? $signed(w_78) : $signed(_GEN_20070); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20667 = 6'h14 == state ? $signed(w_79) : $signed(_GEN_20071); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_20668 = 6'h14 == state ? $signed(temp) : $signed(_GEN_20072); // @[digest.scala 38:19 81:19]
  wire  _GEN_20669 = 6'h14 == state ? 1'h0 : _GEN_20073; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_20672 = 6'h14 == state ? $signed(t) : $signed(_GEN_20076); // @[digest.scala 35:16 81:19]
  wire  _GEN_20673 = 6'h14 == state ? 1'h0 : _GEN_20077; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_20676 = 6'h14 == state ? $signed(e) : $signed(_GEN_20080); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_20677 = 6'h14 == state ? $signed(d) : $signed(_GEN_20081); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_20678 = 6'h14 == state ? $signed(c) : $signed(_GEN_20082); // @[digest.scala 26:16 81:19]
  wire  _GEN_20679 = 6'h14 == state ? 1'h0 : _GEN_20083; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_20682 = 6'h14 == state ? $signed(b) : $signed(_GEN_20086); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_20683 = 6'h14 == state ? $signed(a) : $signed(_GEN_20087); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_20684 = 6'h14 == state ? $signed(i) : $signed(_GEN_20088); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_20766 = 6'h14 == state ? $signed(digest_0) : $signed(_GEN_20170); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20767 = 6'h14 == state ? $signed(digest_1) : $signed(_GEN_20171); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20768 = 6'h14 == state ? $signed(digest_2) : $signed(_GEN_20172); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20769 = 6'h14 == state ? $signed(digest_3) : $signed(_GEN_20173); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20770 = 6'h14 == state ? $signed(digest_4) : $signed(_GEN_20174); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20771 = 6'h14 == state ? $signed(digest_5) : $signed(_GEN_20175); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20772 = 6'h14 == state ? $signed(digest_6) : $signed(_GEN_20176); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20773 = 6'h14 == state ? $signed(digest_7) : $signed(_GEN_20177); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20774 = 6'h14 == state ? $signed(digest_8) : $signed(_GEN_20178); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20775 = 6'h14 == state ? $signed(digest_9) : $signed(_GEN_20179); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20776 = 6'h14 == state ? $signed(digest_10) : $signed(_GEN_20180); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20777 = 6'h14 == state ? $signed(digest_11) : $signed(_GEN_20181); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20778 = 6'h14 == state ? $signed(digest_12) : $signed(_GEN_20182); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20779 = 6'h14 == state ? $signed(digest_13) : $signed(_GEN_20183); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20780 = 6'h14 == state ? $signed(digest_14) : $signed(_GEN_20184); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20781 = 6'h14 == state ? $signed(digest_15) : $signed(_GEN_20185); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20782 = 6'h14 == state ? $signed(digest_16) : $signed(_GEN_20186); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20783 = 6'h14 == state ? $signed(digest_17) : $signed(_GEN_20187); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20784 = 6'h14 == state ? $signed(digest_18) : $signed(_GEN_20188); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20785 = 6'h14 == state ? $signed(digest_19) : $signed(_GEN_20189); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20786 = 6'h14 == state ? $signed(digest_20) : $signed(_GEN_20190); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20787 = 6'h14 == state ? $signed(digest_21) : $signed(_GEN_20191); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20788 = 6'h14 == state ? $signed(digest_22) : $signed(_GEN_20192); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20789 = 6'h14 == state ? $signed(digest_23) : $signed(_GEN_20193); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20790 = 6'h14 == state ? $signed(digest_24) : $signed(_GEN_20194); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20791 = 6'h14 == state ? $signed(digest_25) : $signed(_GEN_20195); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20792 = 6'h14 == state ? $signed(digest_26) : $signed(_GEN_20196); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20793 = 6'h14 == state ? $signed(digest_27) : $signed(_GEN_20197); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20794 = 6'h14 == state ? $signed(digest_28) : $signed(_GEN_20198); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20795 = 6'h14 == state ? $signed(digest_29) : $signed(_GEN_20199); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20796 = 6'h14 == state ? $signed(digest_30) : $signed(_GEN_20200); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20797 = 6'h14 == state ? $signed(digest_31) : $signed(_GEN_20201); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20798 = 6'h14 == state ? $signed(digest_32) : $signed(_GEN_20202); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20799 = 6'h14 == state ? $signed(digest_33) : $signed(_GEN_20203); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20800 = 6'h14 == state ? $signed(digest_34) : $signed(_GEN_20204); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20801 = 6'h14 == state ? $signed(digest_35) : $signed(_GEN_20205); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20802 = 6'h14 == state ? $signed(digest_36) : $signed(_GEN_20206); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20803 = 6'h14 == state ? $signed(digest_37) : $signed(_GEN_20207); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20804 = 6'h14 == state ? $signed(digest_38) : $signed(_GEN_20208); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20805 = 6'h14 == state ? $signed(digest_39) : $signed(_GEN_20209); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20806 = 6'h14 == state ? $signed(digest_40) : $signed(_GEN_20210); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20807 = 6'h14 == state ? $signed(digest_41) : $signed(_GEN_20211); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20808 = 6'h14 == state ? $signed(digest_42) : $signed(_GEN_20212); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20809 = 6'h14 == state ? $signed(digest_43) : $signed(_GEN_20213); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20810 = 6'h14 == state ? $signed(digest_44) : $signed(_GEN_20214); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20811 = 6'h14 == state ? $signed(digest_45) : $signed(_GEN_20215); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20812 = 6'h14 == state ? $signed(digest_46) : $signed(_GEN_20216); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20813 = 6'h14 == state ? $signed(digest_47) : $signed(_GEN_20217); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20814 = 6'h14 == state ? $signed(digest_48) : $signed(_GEN_20218); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20815 = 6'h14 == state ? $signed(digest_49) : $signed(_GEN_20219); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20816 = 6'h14 == state ? $signed(digest_50) : $signed(_GEN_20220); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20817 = 6'h14 == state ? $signed(digest_51) : $signed(_GEN_20221); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20818 = 6'h14 == state ? $signed(digest_52) : $signed(_GEN_20222); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20819 = 6'h14 == state ? $signed(digest_53) : $signed(_GEN_20223); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20820 = 6'h14 == state ? $signed(digest_54) : $signed(_GEN_20224); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20821 = 6'h14 == state ? $signed(digest_55) : $signed(_GEN_20225); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20822 = 6'h14 == state ? $signed(digest_56) : $signed(_GEN_20226); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20823 = 6'h14 == state ? $signed(digest_57) : $signed(_GEN_20227); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20824 = 6'h14 == state ? $signed(digest_58) : $signed(_GEN_20228); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20825 = 6'h14 == state ? $signed(digest_59) : $signed(_GEN_20229); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20826 = 6'h14 == state ? $signed(digest_60) : $signed(_GEN_20230); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20827 = 6'h14 == state ? $signed(digest_61) : $signed(_GEN_20231); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20828 = 6'h14 == state ? $signed(digest_62) : $signed(_GEN_20232); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20829 = 6'h14 == state ? $signed(digest_63) : $signed(_GEN_20233); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20830 = 6'h14 == state ? $signed(digest_64) : $signed(_GEN_20234); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20831 = 6'h14 == state ? $signed(digest_65) : $signed(_GEN_20235); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20832 = 6'h14 == state ? $signed(digest_66) : $signed(_GEN_20236); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20833 = 6'h14 == state ? $signed(digest_67) : $signed(_GEN_20237); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20834 = 6'h14 == state ? $signed(digest_68) : $signed(_GEN_20238); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20835 = 6'h14 == state ? $signed(digest_69) : $signed(_GEN_20239); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20836 = 6'h14 == state ? $signed(digest_70) : $signed(_GEN_20240); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20837 = 6'h14 == state ? $signed(digest_71) : $signed(_GEN_20241); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20838 = 6'h14 == state ? $signed(digest_72) : $signed(_GEN_20242); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20839 = 6'h14 == state ? $signed(digest_73) : $signed(_GEN_20243); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20840 = 6'h14 == state ? $signed(digest_74) : $signed(_GEN_20244); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20841 = 6'h14 == state ? $signed(digest_75) : $signed(_GEN_20245); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20842 = 6'h14 == state ? $signed(digest_76) : $signed(_GEN_20246); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20843 = 6'h14 == state ? $signed(digest_77) : $signed(_GEN_20247); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20844 = 6'h14 == state ? $signed(digest_78) : $signed(_GEN_20248); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_20845 = 6'h14 == state ? $signed(digest_79) : $signed(_GEN_20249); // @[digest.scala 81:19 53:21]
  wire  _GEN_20847 = 6'h14 == state ? 1'h0 : _GEN_20251; // @[digest.scala 81:19 58:25]
  wire  _GEN_20930 = 6'h14 == state ? 1'h0 : _GEN_20334; // @[digest.scala 81:19 63:25]
  wire  _GEN_21013 = 6'h14 == state ? 1'h0 : _GEN_20417; // @[digest.scala 81:19 68:25]
  wire  _GEN_21096 = 6'h14 == state ? 1'h0 : _GEN_20500; // @[digest.scala 81:19 73:25]
  wire  _GEN_21179 = 6'h14 == state ? 1'h0 : _GEN_20583; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_21180 = 6'h13 == state ? $signed(c) : $signed(oldc); // @[digest.scala 160:18 31:19 81:19]
  wire [5:0] _GEN_21181 = 6'h13 == state ? 6'h14 : _GEN_20585; // @[digest.scala 161:19 81:19]
  wire [31:0] _GEN_21182 = 6'h13 == state ? $signed(oldd) : $signed(_GEN_20584); // @[digest.scala 32:19 81:19]
  wire [31:0] _GEN_21183 = 6'h13 == state ? $signed(olde) : $signed(_GEN_20586); // @[digest.scala 33:19 81:19]
  wire [31:0] _GEN_21184 = 6'h13 == state ? $signed(j) : $signed(_GEN_20587); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_21185 = 6'h13 == state ? $signed(w_0) : $signed(_GEN_20588); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21186 = 6'h13 == state ? $signed(w_1) : $signed(_GEN_20589); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21187 = 6'h13 == state ? $signed(w_2) : $signed(_GEN_20590); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21188 = 6'h13 == state ? $signed(w_3) : $signed(_GEN_20591); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21189 = 6'h13 == state ? $signed(w_4) : $signed(_GEN_20592); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21190 = 6'h13 == state ? $signed(w_5) : $signed(_GEN_20593); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21191 = 6'h13 == state ? $signed(w_6) : $signed(_GEN_20594); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21192 = 6'h13 == state ? $signed(w_7) : $signed(_GEN_20595); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21193 = 6'h13 == state ? $signed(w_8) : $signed(_GEN_20596); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21194 = 6'h13 == state ? $signed(w_9) : $signed(_GEN_20597); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21195 = 6'h13 == state ? $signed(w_10) : $signed(_GEN_20598); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21196 = 6'h13 == state ? $signed(w_11) : $signed(_GEN_20599); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21197 = 6'h13 == state ? $signed(w_12) : $signed(_GEN_20600); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21198 = 6'h13 == state ? $signed(w_13) : $signed(_GEN_20601); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21199 = 6'h13 == state ? $signed(w_14) : $signed(_GEN_20602); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21200 = 6'h13 == state ? $signed(w_15) : $signed(_GEN_20603); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21201 = 6'h13 == state ? $signed(w_16) : $signed(_GEN_20604); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21202 = 6'h13 == state ? $signed(w_17) : $signed(_GEN_20605); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21203 = 6'h13 == state ? $signed(w_18) : $signed(_GEN_20606); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21204 = 6'h13 == state ? $signed(w_19) : $signed(_GEN_20607); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21205 = 6'h13 == state ? $signed(w_20) : $signed(_GEN_20608); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21206 = 6'h13 == state ? $signed(w_21) : $signed(_GEN_20609); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21207 = 6'h13 == state ? $signed(w_22) : $signed(_GEN_20610); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21208 = 6'h13 == state ? $signed(w_23) : $signed(_GEN_20611); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21209 = 6'h13 == state ? $signed(w_24) : $signed(_GEN_20612); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21210 = 6'h13 == state ? $signed(w_25) : $signed(_GEN_20613); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21211 = 6'h13 == state ? $signed(w_26) : $signed(_GEN_20614); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21212 = 6'h13 == state ? $signed(w_27) : $signed(_GEN_20615); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21213 = 6'h13 == state ? $signed(w_28) : $signed(_GEN_20616); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21214 = 6'h13 == state ? $signed(w_29) : $signed(_GEN_20617); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21215 = 6'h13 == state ? $signed(w_30) : $signed(_GEN_20618); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21216 = 6'h13 == state ? $signed(w_31) : $signed(_GEN_20619); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21217 = 6'h13 == state ? $signed(w_32) : $signed(_GEN_20620); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21218 = 6'h13 == state ? $signed(w_33) : $signed(_GEN_20621); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21219 = 6'h13 == state ? $signed(w_34) : $signed(_GEN_20622); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21220 = 6'h13 == state ? $signed(w_35) : $signed(_GEN_20623); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21221 = 6'h13 == state ? $signed(w_36) : $signed(_GEN_20624); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21222 = 6'h13 == state ? $signed(w_37) : $signed(_GEN_20625); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21223 = 6'h13 == state ? $signed(w_38) : $signed(_GEN_20626); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21224 = 6'h13 == state ? $signed(w_39) : $signed(_GEN_20627); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21225 = 6'h13 == state ? $signed(w_40) : $signed(_GEN_20628); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21226 = 6'h13 == state ? $signed(w_41) : $signed(_GEN_20629); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21227 = 6'h13 == state ? $signed(w_42) : $signed(_GEN_20630); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21228 = 6'h13 == state ? $signed(w_43) : $signed(_GEN_20631); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21229 = 6'h13 == state ? $signed(w_44) : $signed(_GEN_20632); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21230 = 6'h13 == state ? $signed(w_45) : $signed(_GEN_20633); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21231 = 6'h13 == state ? $signed(w_46) : $signed(_GEN_20634); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21232 = 6'h13 == state ? $signed(w_47) : $signed(_GEN_20635); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21233 = 6'h13 == state ? $signed(w_48) : $signed(_GEN_20636); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21234 = 6'h13 == state ? $signed(w_49) : $signed(_GEN_20637); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21235 = 6'h13 == state ? $signed(w_50) : $signed(_GEN_20638); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21236 = 6'h13 == state ? $signed(w_51) : $signed(_GEN_20639); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21237 = 6'h13 == state ? $signed(w_52) : $signed(_GEN_20640); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21238 = 6'h13 == state ? $signed(w_53) : $signed(_GEN_20641); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21239 = 6'h13 == state ? $signed(w_54) : $signed(_GEN_20642); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21240 = 6'h13 == state ? $signed(w_55) : $signed(_GEN_20643); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21241 = 6'h13 == state ? $signed(w_56) : $signed(_GEN_20644); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21242 = 6'h13 == state ? $signed(w_57) : $signed(_GEN_20645); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21243 = 6'h13 == state ? $signed(w_58) : $signed(_GEN_20646); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21244 = 6'h13 == state ? $signed(w_59) : $signed(_GEN_20647); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21245 = 6'h13 == state ? $signed(w_60) : $signed(_GEN_20648); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21246 = 6'h13 == state ? $signed(w_61) : $signed(_GEN_20649); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21247 = 6'h13 == state ? $signed(w_62) : $signed(_GEN_20650); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21248 = 6'h13 == state ? $signed(w_63) : $signed(_GEN_20651); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21249 = 6'h13 == state ? $signed(w_64) : $signed(_GEN_20652); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21250 = 6'h13 == state ? $signed(w_65) : $signed(_GEN_20653); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21251 = 6'h13 == state ? $signed(w_66) : $signed(_GEN_20654); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21252 = 6'h13 == state ? $signed(w_67) : $signed(_GEN_20655); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21253 = 6'h13 == state ? $signed(w_68) : $signed(_GEN_20656); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21254 = 6'h13 == state ? $signed(w_69) : $signed(_GEN_20657); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21255 = 6'h13 == state ? $signed(w_70) : $signed(_GEN_20658); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21256 = 6'h13 == state ? $signed(w_71) : $signed(_GEN_20659); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21257 = 6'h13 == state ? $signed(w_72) : $signed(_GEN_20660); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21258 = 6'h13 == state ? $signed(w_73) : $signed(_GEN_20661); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21259 = 6'h13 == state ? $signed(w_74) : $signed(_GEN_20662); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21260 = 6'h13 == state ? $signed(w_75) : $signed(_GEN_20663); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21261 = 6'h13 == state ? $signed(w_76) : $signed(_GEN_20664); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21262 = 6'h13 == state ? $signed(w_77) : $signed(_GEN_20665); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21263 = 6'h13 == state ? $signed(w_78) : $signed(_GEN_20666); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21264 = 6'h13 == state ? $signed(w_79) : $signed(_GEN_20667); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21265 = 6'h13 == state ? $signed(temp) : $signed(_GEN_20668); // @[digest.scala 38:19 81:19]
  wire  _GEN_21266 = 6'h13 == state ? 1'h0 : _GEN_20669; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_21269 = 6'h13 == state ? $signed(t) : $signed(_GEN_20672); // @[digest.scala 35:16 81:19]
  wire  _GEN_21270 = 6'h13 == state ? 1'h0 : _GEN_20673; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_21273 = 6'h13 == state ? $signed(e) : $signed(_GEN_20676); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_21274 = 6'h13 == state ? $signed(d) : $signed(_GEN_20677); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_21275 = 6'h13 == state ? $signed(c) : $signed(_GEN_20678); // @[digest.scala 26:16 81:19]
  wire  _GEN_21276 = 6'h13 == state ? 1'h0 : _GEN_20679; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_21279 = 6'h13 == state ? $signed(b) : $signed(_GEN_20682); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_21280 = 6'h13 == state ? $signed(a) : $signed(_GEN_20683); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_21281 = 6'h13 == state ? $signed(i) : $signed(_GEN_20684); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_21363 = 6'h13 == state ? $signed(digest_0) : $signed(_GEN_20766); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21364 = 6'h13 == state ? $signed(digest_1) : $signed(_GEN_20767); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21365 = 6'h13 == state ? $signed(digest_2) : $signed(_GEN_20768); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21366 = 6'h13 == state ? $signed(digest_3) : $signed(_GEN_20769); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21367 = 6'h13 == state ? $signed(digest_4) : $signed(_GEN_20770); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21368 = 6'h13 == state ? $signed(digest_5) : $signed(_GEN_20771); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21369 = 6'h13 == state ? $signed(digest_6) : $signed(_GEN_20772); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21370 = 6'h13 == state ? $signed(digest_7) : $signed(_GEN_20773); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21371 = 6'h13 == state ? $signed(digest_8) : $signed(_GEN_20774); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21372 = 6'h13 == state ? $signed(digest_9) : $signed(_GEN_20775); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21373 = 6'h13 == state ? $signed(digest_10) : $signed(_GEN_20776); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21374 = 6'h13 == state ? $signed(digest_11) : $signed(_GEN_20777); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21375 = 6'h13 == state ? $signed(digest_12) : $signed(_GEN_20778); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21376 = 6'h13 == state ? $signed(digest_13) : $signed(_GEN_20779); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21377 = 6'h13 == state ? $signed(digest_14) : $signed(_GEN_20780); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21378 = 6'h13 == state ? $signed(digest_15) : $signed(_GEN_20781); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21379 = 6'h13 == state ? $signed(digest_16) : $signed(_GEN_20782); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21380 = 6'h13 == state ? $signed(digest_17) : $signed(_GEN_20783); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21381 = 6'h13 == state ? $signed(digest_18) : $signed(_GEN_20784); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21382 = 6'h13 == state ? $signed(digest_19) : $signed(_GEN_20785); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21383 = 6'h13 == state ? $signed(digest_20) : $signed(_GEN_20786); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21384 = 6'h13 == state ? $signed(digest_21) : $signed(_GEN_20787); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21385 = 6'h13 == state ? $signed(digest_22) : $signed(_GEN_20788); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21386 = 6'h13 == state ? $signed(digest_23) : $signed(_GEN_20789); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21387 = 6'h13 == state ? $signed(digest_24) : $signed(_GEN_20790); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21388 = 6'h13 == state ? $signed(digest_25) : $signed(_GEN_20791); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21389 = 6'h13 == state ? $signed(digest_26) : $signed(_GEN_20792); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21390 = 6'h13 == state ? $signed(digest_27) : $signed(_GEN_20793); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21391 = 6'h13 == state ? $signed(digest_28) : $signed(_GEN_20794); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21392 = 6'h13 == state ? $signed(digest_29) : $signed(_GEN_20795); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21393 = 6'h13 == state ? $signed(digest_30) : $signed(_GEN_20796); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21394 = 6'h13 == state ? $signed(digest_31) : $signed(_GEN_20797); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21395 = 6'h13 == state ? $signed(digest_32) : $signed(_GEN_20798); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21396 = 6'h13 == state ? $signed(digest_33) : $signed(_GEN_20799); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21397 = 6'h13 == state ? $signed(digest_34) : $signed(_GEN_20800); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21398 = 6'h13 == state ? $signed(digest_35) : $signed(_GEN_20801); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21399 = 6'h13 == state ? $signed(digest_36) : $signed(_GEN_20802); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21400 = 6'h13 == state ? $signed(digest_37) : $signed(_GEN_20803); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21401 = 6'h13 == state ? $signed(digest_38) : $signed(_GEN_20804); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21402 = 6'h13 == state ? $signed(digest_39) : $signed(_GEN_20805); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21403 = 6'h13 == state ? $signed(digest_40) : $signed(_GEN_20806); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21404 = 6'h13 == state ? $signed(digest_41) : $signed(_GEN_20807); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21405 = 6'h13 == state ? $signed(digest_42) : $signed(_GEN_20808); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21406 = 6'h13 == state ? $signed(digest_43) : $signed(_GEN_20809); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21407 = 6'h13 == state ? $signed(digest_44) : $signed(_GEN_20810); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21408 = 6'h13 == state ? $signed(digest_45) : $signed(_GEN_20811); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21409 = 6'h13 == state ? $signed(digest_46) : $signed(_GEN_20812); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21410 = 6'h13 == state ? $signed(digest_47) : $signed(_GEN_20813); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21411 = 6'h13 == state ? $signed(digest_48) : $signed(_GEN_20814); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21412 = 6'h13 == state ? $signed(digest_49) : $signed(_GEN_20815); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21413 = 6'h13 == state ? $signed(digest_50) : $signed(_GEN_20816); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21414 = 6'h13 == state ? $signed(digest_51) : $signed(_GEN_20817); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21415 = 6'h13 == state ? $signed(digest_52) : $signed(_GEN_20818); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21416 = 6'h13 == state ? $signed(digest_53) : $signed(_GEN_20819); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21417 = 6'h13 == state ? $signed(digest_54) : $signed(_GEN_20820); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21418 = 6'h13 == state ? $signed(digest_55) : $signed(_GEN_20821); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21419 = 6'h13 == state ? $signed(digest_56) : $signed(_GEN_20822); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21420 = 6'h13 == state ? $signed(digest_57) : $signed(_GEN_20823); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21421 = 6'h13 == state ? $signed(digest_58) : $signed(_GEN_20824); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21422 = 6'h13 == state ? $signed(digest_59) : $signed(_GEN_20825); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21423 = 6'h13 == state ? $signed(digest_60) : $signed(_GEN_20826); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21424 = 6'h13 == state ? $signed(digest_61) : $signed(_GEN_20827); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21425 = 6'h13 == state ? $signed(digest_62) : $signed(_GEN_20828); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21426 = 6'h13 == state ? $signed(digest_63) : $signed(_GEN_20829); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21427 = 6'h13 == state ? $signed(digest_64) : $signed(_GEN_20830); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21428 = 6'h13 == state ? $signed(digest_65) : $signed(_GEN_20831); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21429 = 6'h13 == state ? $signed(digest_66) : $signed(_GEN_20832); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21430 = 6'h13 == state ? $signed(digest_67) : $signed(_GEN_20833); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21431 = 6'h13 == state ? $signed(digest_68) : $signed(_GEN_20834); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21432 = 6'h13 == state ? $signed(digest_69) : $signed(_GEN_20835); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21433 = 6'h13 == state ? $signed(digest_70) : $signed(_GEN_20836); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21434 = 6'h13 == state ? $signed(digest_71) : $signed(_GEN_20837); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21435 = 6'h13 == state ? $signed(digest_72) : $signed(_GEN_20838); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21436 = 6'h13 == state ? $signed(digest_73) : $signed(_GEN_20839); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21437 = 6'h13 == state ? $signed(digest_74) : $signed(_GEN_20840); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21438 = 6'h13 == state ? $signed(digest_75) : $signed(_GEN_20841); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21439 = 6'h13 == state ? $signed(digest_76) : $signed(_GEN_20842); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21440 = 6'h13 == state ? $signed(digest_77) : $signed(_GEN_20843); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21441 = 6'h13 == state ? $signed(digest_78) : $signed(_GEN_20844); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21442 = 6'h13 == state ? $signed(digest_79) : $signed(_GEN_20845); // @[digest.scala 81:19 53:21]
  wire  _GEN_21444 = 6'h13 == state ? 1'h0 : _GEN_20847; // @[digest.scala 81:19 58:25]
  wire  _GEN_21527 = 6'h13 == state ? 1'h0 : _GEN_20930; // @[digest.scala 81:19 63:25]
  wire  _GEN_21610 = 6'h13 == state ? 1'h0 : _GEN_21013; // @[digest.scala 81:19 68:25]
  wire  _GEN_21693 = 6'h13 == state ? 1'h0 : _GEN_21096; // @[digest.scala 81:19 73:25]
  wire  _GEN_21776 = 6'h13 == state ? 1'h0 : _GEN_21179; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_21777 = 6'h12 == state ? $signed(b) : $signed(oldb); // @[digest.scala 156:18 30:19 81:19]
  wire [5:0] _GEN_21778 = 6'h12 == state ? 6'h13 : _GEN_21181; // @[digest.scala 157:19 81:19]
  wire [31:0] _GEN_21779 = 6'h12 == state ? $signed(oldc) : $signed(_GEN_21180); // @[digest.scala 31:19 81:19]
  wire [31:0] _GEN_21780 = 6'h12 == state ? $signed(oldd) : $signed(_GEN_21182); // @[digest.scala 32:19 81:19]
  wire [31:0] _GEN_21781 = 6'h12 == state ? $signed(olde) : $signed(_GEN_21183); // @[digest.scala 33:19 81:19]
  wire [31:0] _GEN_21782 = 6'h12 == state ? $signed(j) : $signed(_GEN_21184); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_21783 = 6'h12 == state ? $signed(w_0) : $signed(_GEN_21185); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21784 = 6'h12 == state ? $signed(w_1) : $signed(_GEN_21186); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21785 = 6'h12 == state ? $signed(w_2) : $signed(_GEN_21187); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21786 = 6'h12 == state ? $signed(w_3) : $signed(_GEN_21188); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21787 = 6'h12 == state ? $signed(w_4) : $signed(_GEN_21189); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21788 = 6'h12 == state ? $signed(w_5) : $signed(_GEN_21190); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21789 = 6'h12 == state ? $signed(w_6) : $signed(_GEN_21191); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21790 = 6'h12 == state ? $signed(w_7) : $signed(_GEN_21192); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21791 = 6'h12 == state ? $signed(w_8) : $signed(_GEN_21193); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21792 = 6'h12 == state ? $signed(w_9) : $signed(_GEN_21194); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21793 = 6'h12 == state ? $signed(w_10) : $signed(_GEN_21195); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21794 = 6'h12 == state ? $signed(w_11) : $signed(_GEN_21196); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21795 = 6'h12 == state ? $signed(w_12) : $signed(_GEN_21197); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21796 = 6'h12 == state ? $signed(w_13) : $signed(_GEN_21198); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21797 = 6'h12 == state ? $signed(w_14) : $signed(_GEN_21199); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21798 = 6'h12 == state ? $signed(w_15) : $signed(_GEN_21200); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21799 = 6'h12 == state ? $signed(w_16) : $signed(_GEN_21201); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21800 = 6'h12 == state ? $signed(w_17) : $signed(_GEN_21202); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21801 = 6'h12 == state ? $signed(w_18) : $signed(_GEN_21203); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21802 = 6'h12 == state ? $signed(w_19) : $signed(_GEN_21204); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21803 = 6'h12 == state ? $signed(w_20) : $signed(_GEN_21205); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21804 = 6'h12 == state ? $signed(w_21) : $signed(_GEN_21206); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21805 = 6'h12 == state ? $signed(w_22) : $signed(_GEN_21207); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21806 = 6'h12 == state ? $signed(w_23) : $signed(_GEN_21208); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21807 = 6'h12 == state ? $signed(w_24) : $signed(_GEN_21209); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21808 = 6'h12 == state ? $signed(w_25) : $signed(_GEN_21210); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21809 = 6'h12 == state ? $signed(w_26) : $signed(_GEN_21211); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21810 = 6'h12 == state ? $signed(w_27) : $signed(_GEN_21212); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21811 = 6'h12 == state ? $signed(w_28) : $signed(_GEN_21213); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21812 = 6'h12 == state ? $signed(w_29) : $signed(_GEN_21214); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21813 = 6'h12 == state ? $signed(w_30) : $signed(_GEN_21215); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21814 = 6'h12 == state ? $signed(w_31) : $signed(_GEN_21216); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21815 = 6'h12 == state ? $signed(w_32) : $signed(_GEN_21217); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21816 = 6'h12 == state ? $signed(w_33) : $signed(_GEN_21218); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21817 = 6'h12 == state ? $signed(w_34) : $signed(_GEN_21219); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21818 = 6'h12 == state ? $signed(w_35) : $signed(_GEN_21220); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21819 = 6'h12 == state ? $signed(w_36) : $signed(_GEN_21221); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21820 = 6'h12 == state ? $signed(w_37) : $signed(_GEN_21222); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21821 = 6'h12 == state ? $signed(w_38) : $signed(_GEN_21223); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21822 = 6'h12 == state ? $signed(w_39) : $signed(_GEN_21224); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21823 = 6'h12 == state ? $signed(w_40) : $signed(_GEN_21225); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21824 = 6'h12 == state ? $signed(w_41) : $signed(_GEN_21226); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21825 = 6'h12 == state ? $signed(w_42) : $signed(_GEN_21227); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21826 = 6'h12 == state ? $signed(w_43) : $signed(_GEN_21228); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21827 = 6'h12 == state ? $signed(w_44) : $signed(_GEN_21229); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21828 = 6'h12 == state ? $signed(w_45) : $signed(_GEN_21230); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21829 = 6'h12 == state ? $signed(w_46) : $signed(_GEN_21231); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21830 = 6'h12 == state ? $signed(w_47) : $signed(_GEN_21232); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21831 = 6'h12 == state ? $signed(w_48) : $signed(_GEN_21233); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21832 = 6'h12 == state ? $signed(w_49) : $signed(_GEN_21234); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21833 = 6'h12 == state ? $signed(w_50) : $signed(_GEN_21235); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21834 = 6'h12 == state ? $signed(w_51) : $signed(_GEN_21236); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21835 = 6'h12 == state ? $signed(w_52) : $signed(_GEN_21237); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21836 = 6'h12 == state ? $signed(w_53) : $signed(_GEN_21238); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21837 = 6'h12 == state ? $signed(w_54) : $signed(_GEN_21239); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21838 = 6'h12 == state ? $signed(w_55) : $signed(_GEN_21240); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21839 = 6'h12 == state ? $signed(w_56) : $signed(_GEN_21241); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21840 = 6'h12 == state ? $signed(w_57) : $signed(_GEN_21242); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21841 = 6'h12 == state ? $signed(w_58) : $signed(_GEN_21243); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21842 = 6'h12 == state ? $signed(w_59) : $signed(_GEN_21244); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21843 = 6'h12 == state ? $signed(w_60) : $signed(_GEN_21245); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21844 = 6'h12 == state ? $signed(w_61) : $signed(_GEN_21246); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21845 = 6'h12 == state ? $signed(w_62) : $signed(_GEN_21247); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21846 = 6'h12 == state ? $signed(w_63) : $signed(_GEN_21248); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21847 = 6'h12 == state ? $signed(w_64) : $signed(_GEN_21249); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21848 = 6'h12 == state ? $signed(w_65) : $signed(_GEN_21250); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21849 = 6'h12 == state ? $signed(w_66) : $signed(_GEN_21251); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21850 = 6'h12 == state ? $signed(w_67) : $signed(_GEN_21252); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21851 = 6'h12 == state ? $signed(w_68) : $signed(_GEN_21253); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21852 = 6'h12 == state ? $signed(w_69) : $signed(_GEN_21254); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21853 = 6'h12 == state ? $signed(w_70) : $signed(_GEN_21255); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21854 = 6'h12 == state ? $signed(w_71) : $signed(_GEN_21256); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21855 = 6'h12 == state ? $signed(w_72) : $signed(_GEN_21257); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21856 = 6'h12 == state ? $signed(w_73) : $signed(_GEN_21258); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21857 = 6'h12 == state ? $signed(w_74) : $signed(_GEN_21259); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21858 = 6'h12 == state ? $signed(w_75) : $signed(_GEN_21260); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21859 = 6'h12 == state ? $signed(w_76) : $signed(_GEN_21261); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21860 = 6'h12 == state ? $signed(w_77) : $signed(_GEN_21262); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21861 = 6'h12 == state ? $signed(w_78) : $signed(_GEN_21263); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21862 = 6'h12 == state ? $signed(w_79) : $signed(_GEN_21264); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_21863 = 6'h12 == state ? $signed(temp) : $signed(_GEN_21265); // @[digest.scala 38:19 81:19]
  wire  _GEN_21864 = 6'h12 == state ? 1'h0 : _GEN_21266; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_21867 = 6'h12 == state ? $signed(t) : $signed(_GEN_21269); // @[digest.scala 35:16 81:19]
  wire  _GEN_21868 = 6'h12 == state ? 1'h0 : _GEN_21270; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_21871 = 6'h12 == state ? $signed(e) : $signed(_GEN_21273); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_21872 = 6'h12 == state ? $signed(d) : $signed(_GEN_21274); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_21873 = 6'h12 == state ? $signed(c) : $signed(_GEN_21275); // @[digest.scala 26:16 81:19]
  wire  _GEN_21874 = 6'h12 == state ? 1'h0 : _GEN_21276; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_21877 = 6'h12 == state ? $signed(b) : $signed(_GEN_21279); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_21878 = 6'h12 == state ? $signed(a) : $signed(_GEN_21280); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_21879 = 6'h12 == state ? $signed(i) : $signed(_GEN_21281); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_21961 = 6'h12 == state ? $signed(digest_0) : $signed(_GEN_21363); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21962 = 6'h12 == state ? $signed(digest_1) : $signed(_GEN_21364); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21963 = 6'h12 == state ? $signed(digest_2) : $signed(_GEN_21365); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21964 = 6'h12 == state ? $signed(digest_3) : $signed(_GEN_21366); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21965 = 6'h12 == state ? $signed(digest_4) : $signed(_GEN_21367); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21966 = 6'h12 == state ? $signed(digest_5) : $signed(_GEN_21368); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21967 = 6'h12 == state ? $signed(digest_6) : $signed(_GEN_21369); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21968 = 6'h12 == state ? $signed(digest_7) : $signed(_GEN_21370); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21969 = 6'h12 == state ? $signed(digest_8) : $signed(_GEN_21371); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21970 = 6'h12 == state ? $signed(digest_9) : $signed(_GEN_21372); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21971 = 6'h12 == state ? $signed(digest_10) : $signed(_GEN_21373); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21972 = 6'h12 == state ? $signed(digest_11) : $signed(_GEN_21374); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21973 = 6'h12 == state ? $signed(digest_12) : $signed(_GEN_21375); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21974 = 6'h12 == state ? $signed(digest_13) : $signed(_GEN_21376); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21975 = 6'h12 == state ? $signed(digest_14) : $signed(_GEN_21377); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21976 = 6'h12 == state ? $signed(digest_15) : $signed(_GEN_21378); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21977 = 6'h12 == state ? $signed(digest_16) : $signed(_GEN_21379); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21978 = 6'h12 == state ? $signed(digest_17) : $signed(_GEN_21380); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21979 = 6'h12 == state ? $signed(digest_18) : $signed(_GEN_21381); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21980 = 6'h12 == state ? $signed(digest_19) : $signed(_GEN_21382); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21981 = 6'h12 == state ? $signed(digest_20) : $signed(_GEN_21383); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21982 = 6'h12 == state ? $signed(digest_21) : $signed(_GEN_21384); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21983 = 6'h12 == state ? $signed(digest_22) : $signed(_GEN_21385); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21984 = 6'h12 == state ? $signed(digest_23) : $signed(_GEN_21386); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21985 = 6'h12 == state ? $signed(digest_24) : $signed(_GEN_21387); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21986 = 6'h12 == state ? $signed(digest_25) : $signed(_GEN_21388); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21987 = 6'h12 == state ? $signed(digest_26) : $signed(_GEN_21389); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21988 = 6'h12 == state ? $signed(digest_27) : $signed(_GEN_21390); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21989 = 6'h12 == state ? $signed(digest_28) : $signed(_GEN_21391); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21990 = 6'h12 == state ? $signed(digest_29) : $signed(_GEN_21392); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21991 = 6'h12 == state ? $signed(digest_30) : $signed(_GEN_21393); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21992 = 6'h12 == state ? $signed(digest_31) : $signed(_GEN_21394); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21993 = 6'h12 == state ? $signed(digest_32) : $signed(_GEN_21395); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21994 = 6'h12 == state ? $signed(digest_33) : $signed(_GEN_21396); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21995 = 6'h12 == state ? $signed(digest_34) : $signed(_GEN_21397); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21996 = 6'h12 == state ? $signed(digest_35) : $signed(_GEN_21398); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21997 = 6'h12 == state ? $signed(digest_36) : $signed(_GEN_21399); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21998 = 6'h12 == state ? $signed(digest_37) : $signed(_GEN_21400); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_21999 = 6'h12 == state ? $signed(digest_38) : $signed(_GEN_21401); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22000 = 6'h12 == state ? $signed(digest_39) : $signed(_GEN_21402); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22001 = 6'h12 == state ? $signed(digest_40) : $signed(_GEN_21403); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22002 = 6'h12 == state ? $signed(digest_41) : $signed(_GEN_21404); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22003 = 6'h12 == state ? $signed(digest_42) : $signed(_GEN_21405); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22004 = 6'h12 == state ? $signed(digest_43) : $signed(_GEN_21406); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22005 = 6'h12 == state ? $signed(digest_44) : $signed(_GEN_21407); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22006 = 6'h12 == state ? $signed(digest_45) : $signed(_GEN_21408); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22007 = 6'h12 == state ? $signed(digest_46) : $signed(_GEN_21409); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22008 = 6'h12 == state ? $signed(digest_47) : $signed(_GEN_21410); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22009 = 6'h12 == state ? $signed(digest_48) : $signed(_GEN_21411); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22010 = 6'h12 == state ? $signed(digest_49) : $signed(_GEN_21412); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22011 = 6'h12 == state ? $signed(digest_50) : $signed(_GEN_21413); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22012 = 6'h12 == state ? $signed(digest_51) : $signed(_GEN_21414); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22013 = 6'h12 == state ? $signed(digest_52) : $signed(_GEN_21415); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22014 = 6'h12 == state ? $signed(digest_53) : $signed(_GEN_21416); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22015 = 6'h12 == state ? $signed(digest_54) : $signed(_GEN_21417); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22016 = 6'h12 == state ? $signed(digest_55) : $signed(_GEN_21418); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22017 = 6'h12 == state ? $signed(digest_56) : $signed(_GEN_21419); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22018 = 6'h12 == state ? $signed(digest_57) : $signed(_GEN_21420); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22019 = 6'h12 == state ? $signed(digest_58) : $signed(_GEN_21421); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22020 = 6'h12 == state ? $signed(digest_59) : $signed(_GEN_21422); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22021 = 6'h12 == state ? $signed(digest_60) : $signed(_GEN_21423); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22022 = 6'h12 == state ? $signed(digest_61) : $signed(_GEN_21424); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22023 = 6'h12 == state ? $signed(digest_62) : $signed(_GEN_21425); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22024 = 6'h12 == state ? $signed(digest_63) : $signed(_GEN_21426); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22025 = 6'h12 == state ? $signed(digest_64) : $signed(_GEN_21427); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22026 = 6'h12 == state ? $signed(digest_65) : $signed(_GEN_21428); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22027 = 6'h12 == state ? $signed(digest_66) : $signed(_GEN_21429); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22028 = 6'h12 == state ? $signed(digest_67) : $signed(_GEN_21430); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22029 = 6'h12 == state ? $signed(digest_68) : $signed(_GEN_21431); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22030 = 6'h12 == state ? $signed(digest_69) : $signed(_GEN_21432); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22031 = 6'h12 == state ? $signed(digest_70) : $signed(_GEN_21433); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22032 = 6'h12 == state ? $signed(digest_71) : $signed(_GEN_21434); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22033 = 6'h12 == state ? $signed(digest_72) : $signed(_GEN_21435); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22034 = 6'h12 == state ? $signed(digest_73) : $signed(_GEN_21436); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22035 = 6'h12 == state ? $signed(digest_74) : $signed(_GEN_21437); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22036 = 6'h12 == state ? $signed(digest_75) : $signed(_GEN_21438); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22037 = 6'h12 == state ? $signed(digest_76) : $signed(_GEN_21439); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22038 = 6'h12 == state ? $signed(digest_77) : $signed(_GEN_21440); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22039 = 6'h12 == state ? $signed(digest_78) : $signed(_GEN_21441); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22040 = 6'h12 == state ? $signed(digest_79) : $signed(_GEN_21442); // @[digest.scala 81:19 53:21]
  wire  _GEN_22042 = 6'h12 == state ? 1'h0 : _GEN_21444; // @[digest.scala 81:19 58:25]
  wire  _GEN_22125 = 6'h12 == state ? 1'h0 : _GEN_21527; // @[digest.scala 81:19 63:25]
  wire  _GEN_22208 = 6'h12 == state ? 1'h0 : _GEN_21610; // @[digest.scala 81:19 68:25]
  wire  _GEN_22291 = 6'h12 == state ? 1'h0 : _GEN_21693; // @[digest.scala 81:19 73:25]
  wire  _GEN_22374 = 6'h12 == state ? 1'h0 : _GEN_21776; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_22375 = 6'h11 == state ? $signed(a) : $signed(olda); // @[digest.scala 152:18 29:19 81:19]
  wire [5:0] _GEN_22376 = 6'h11 == state ? 6'h12 : _GEN_21778; // @[digest.scala 153:19 81:19]
  wire [31:0] _GEN_22377 = 6'h11 == state ? $signed(oldb) : $signed(_GEN_21777); // @[digest.scala 30:19 81:19]
  wire [31:0] _GEN_22378 = 6'h11 == state ? $signed(oldc) : $signed(_GEN_21779); // @[digest.scala 31:19 81:19]
  wire [31:0] _GEN_22379 = 6'h11 == state ? $signed(oldd) : $signed(_GEN_21780); // @[digest.scala 32:19 81:19]
  wire [31:0] _GEN_22380 = 6'h11 == state ? $signed(olde) : $signed(_GEN_21781); // @[digest.scala 33:19 81:19]
  wire [31:0] _GEN_22381 = 6'h11 == state ? $signed(j) : $signed(_GEN_21782); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_22382 = 6'h11 == state ? $signed(w_0) : $signed(_GEN_21783); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22383 = 6'h11 == state ? $signed(w_1) : $signed(_GEN_21784); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22384 = 6'h11 == state ? $signed(w_2) : $signed(_GEN_21785); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22385 = 6'h11 == state ? $signed(w_3) : $signed(_GEN_21786); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22386 = 6'h11 == state ? $signed(w_4) : $signed(_GEN_21787); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22387 = 6'h11 == state ? $signed(w_5) : $signed(_GEN_21788); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22388 = 6'h11 == state ? $signed(w_6) : $signed(_GEN_21789); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22389 = 6'h11 == state ? $signed(w_7) : $signed(_GEN_21790); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22390 = 6'h11 == state ? $signed(w_8) : $signed(_GEN_21791); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22391 = 6'h11 == state ? $signed(w_9) : $signed(_GEN_21792); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22392 = 6'h11 == state ? $signed(w_10) : $signed(_GEN_21793); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22393 = 6'h11 == state ? $signed(w_11) : $signed(_GEN_21794); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22394 = 6'h11 == state ? $signed(w_12) : $signed(_GEN_21795); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22395 = 6'h11 == state ? $signed(w_13) : $signed(_GEN_21796); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22396 = 6'h11 == state ? $signed(w_14) : $signed(_GEN_21797); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22397 = 6'h11 == state ? $signed(w_15) : $signed(_GEN_21798); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22398 = 6'h11 == state ? $signed(w_16) : $signed(_GEN_21799); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22399 = 6'h11 == state ? $signed(w_17) : $signed(_GEN_21800); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22400 = 6'h11 == state ? $signed(w_18) : $signed(_GEN_21801); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22401 = 6'h11 == state ? $signed(w_19) : $signed(_GEN_21802); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22402 = 6'h11 == state ? $signed(w_20) : $signed(_GEN_21803); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22403 = 6'h11 == state ? $signed(w_21) : $signed(_GEN_21804); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22404 = 6'h11 == state ? $signed(w_22) : $signed(_GEN_21805); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22405 = 6'h11 == state ? $signed(w_23) : $signed(_GEN_21806); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22406 = 6'h11 == state ? $signed(w_24) : $signed(_GEN_21807); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22407 = 6'h11 == state ? $signed(w_25) : $signed(_GEN_21808); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22408 = 6'h11 == state ? $signed(w_26) : $signed(_GEN_21809); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22409 = 6'h11 == state ? $signed(w_27) : $signed(_GEN_21810); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22410 = 6'h11 == state ? $signed(w_28) : $signed(_GEN_21811); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22411 = 6'h11 == state ? $signed(w_29) : $signed(_GEN_21812); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22412 = 6'h11 == state ? $signed(w_30) : $signed(_GEN_21813); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22413 = 6'h11 == state ? $signed(w_31) : $signed(_GEN_21814); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22414 = 6'h11 == state ? $signed(w_32) : $signed(_GEN_21815); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22415 = 6'h11 == state ? $signed(w_33) : $signed(_GEN_21816); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22416 = 6'h11 == state ? $signed(w_34) : $signed(_GEN_21817); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22417 = 6'h11 == state ? $signed(w_35) : $signed(_GEN_21818); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22418 = 6'h11 == state ? $signed(w_36) : $signed(_GEN_21819); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22419 = 6'h11 == state ? $signed(w_37) : $signed(_GEN_21820); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22420 = 6'h11 == state ? $signed(w_38) : $signed(_GEN_21821); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22421 = 6'h11 == state ? $signed(w_39) : $signed(_GEN_21822); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22422 = 6'h11 == state ? $signed(w_40) : $signed(_GEN_21823); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22423 = 6'h11 == state ? $signed(w_41) : $signed(_GEN_21824); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22424 = 6'h11 == state ? $signed(w_42) : $signed(_GEN_21825); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22425 = 6'h11 == state ? $signed(w_43) : $signed(_GEN_21826); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22426 = 6'h11 == state ? $signed(w_44) : $signed(_GEN_21827); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22427 = 6'h11 == state ? $signed(w_45) : $signed(_GEN_21828); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22428 = 6'h11 == state ? $signed(w_46) : $signed(_GEN_21829); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22429 = 6'h11 == state ? $signed(w_47) : $signed(_GEN_21830); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22430 = 6'h11 == state ? $signed(w_48) : $signed(_GEN_21831); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22431 = 6'h11 == state ? $signed(w_49) : $signed(_GEN_21832); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22432 = 6'h11 == state ? $signed(w_50) : $signed(_GEN_21833); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22433 = 6'h11 == state ? $signed(w_51) : $signed(_GEN_21834); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22434 = 6'h11 == state ? $signed(w_52) : $signed(_GEN_21835); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22435 = 6'h11 == state ? $signed(w_53) : $signed(_GEN_21836); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22436 = 6'h11 == state ? $signed(w_54) : $signed(_GEN_21837); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22437 = 6'h11 == state ? $signed(w_55) : $signed(_GEN_21838); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22438 = 6'h11 == state ? $signed(w_56) : $signed(_GEN_21839); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22439 = 6'h11 == state ? $signed(w_57) : $signed(_GEN_21840); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22440 = 6'h11 == state ? $signed(w_58) : $signed(_GEN_21841); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22441 = 6'h11 == state ? $signed(w_59) : $signed(_GEN_21842); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22442 = 6'h11 == state ? $signed(w_60) : $signed(_GEN_21843); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22443 = 6'h11 == state ? $signed(w_61) : $signed(_GEN_21844); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22444 = 6'h11 == state ? $signed(w_62) : $signed(_GEN_21845); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22445 = 6'h11 == state ? $signed(w_63) : $signed(_GEN_21846); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22446 = 6'h11 == state ? $signed(w_64) : $signed(_GEN_21847); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22447 = 6'h11 == state ? $signed(w_65) : $signed(_GEN_21848); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22448 = 6'h11 == state ? $signed(w_66) : $signed(_GEN_21849); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22449 = 6'h11 == state ? $signed(w_67) : $signed(_GEN_21850); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22450 = 6'h11 == state ? $signed(w_68) : $signed(_GEN_21851); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22451 = 6'h11 == state ? $signed(w_69) : $signed(_GEN_21852); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22452 = 6'h11 == state ? $signed(w_70) : $signed(_GEN_21853); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22453 = 6'h11 == state ? $signed(w_71) : $signed(_GEN_21854); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22454 = 6'h11 == state ? $signed(w_72) : $signed(_GEN_21855); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22455 = 6'h11 == state ? $signed(w_73) : $signed(_GEN_21856); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22456 = 6'h11 == state ? $signed(w_74) : $signed(_GEN_21857); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22457 = 6'h11 == state ? $signed(w_75) : $signed(_GEN_21858); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22458 = 6'h11 == state ? $signed(w_76) : $signed(_GEN_21859); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22459 = 6'h11 == state ? $signed(w_77) : $signed(_GEN_21860); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22460 = 6'h11 == state ? $signed(w_78) : $signed(_GEN_21861); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22461 = 6'h11 == state ? $signed(w_79) : $signed(_GEN_21862); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22462 = 6'h11 == state ? $signed(temp) : $signed(_GEN_21863); // @[digest.scala 38:19 81:19]
  wire  _GEN_22463 = 6'h11 == state ? 1'h0 : _GEN_21864; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_22466 = 6'h11 == state ? $signed(t) : $signed(_GEN_21867); // @[digest.scala 35:16 81:19]
  wire  _GEN_22467 = 6'h11 == state ? 1'h0 : _GEN_21868; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_22470 = 6'h11 == state ? $signed(e) : $signed(_GEN_21871); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_22471 = 6'h11 == state ? $signed(d) : $signed(_GEN_21872); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_22472 = 6'h11 == state ? $signed(c) : $signed(_GEN_21873); // @[digest.scala 26:16 81:19]
  wire  _GEN_22473 = 6'h11 == state ? 1'h0 : _GEN_21874; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_22476 = 6'h11 == state ? $signed(b) : $signed(_GEN_21877); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_22477 = 6'h11 == state ? $signed(a) : $signed(_GEN_21878); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_22478 = 6'h11 == state ? $signed(i) : $signed(_GEN_21879); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_22560 = 6'h11 == state ? $signed(digest_0) : $signed(_GEN_21961); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22561 = 6'h11 == state ? $signed(digest_1) : $signed(_GEN_21962); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22562 = 6'h11 == state ? $signed(digest_2) : $signed(_GEN_21963); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22563 = 6'h11 == state ? $signed(digest_3) : $signed(_GEN_21964); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22564 = 6'h11 == state ? $signed(digest_4) : $signed(_GEN_21965); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22565 = 6'h11 == state ? $signed(digest_5) : $signed(_GEN_21966); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22566 = 6'h11 == state ? $signed(digest_6) : $signed(_GEN_21967); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22567 = 6'h11 == state ? $signed(digest_7) : $signed(_GEN_21968); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22568 = 6'h11 == state ? $signed(digest_8) : $signed(_GEN_21969); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22569 = 6'h11 == state ? $signed(digest_9) : $signed(_GEN_21970); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22570 = 6'h11 == state ? $signed(digest_10) : $signed(_GEN_21971); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22571 = 6'h11 == state ? $signed(digest_11) : $signed(_GEN_21972); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22572 = 6'h11 == state ? $signed(digest_12) : $signed(_GEN_21973); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22573 = 6'h11 == state ? $signed(digest_13) : $signed(_GEN_21974); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22574 = 6'h11 == state ? $signed(digest_14) : $signed(_GEN_21975); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22575 = 6'h11 == state ? $signed(digest_15) : $signed(_GEN_21976); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22576 = 6'h11 == state ? $signed(digest_16) : $signed(_GEN_21977); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22577 = 6'h11 == state ? $signed(digest_17) : $signed(_GEN_21978); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22578 = 6'h11 == state ? $signed(digest_18) : $signed(_GEN_21979); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22579 = 6'h11 == state ? $signed(digest_19) : $signed(_GEN_21980); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22580 = 6'h11 == state ? $signed(digest_20) : $signed(_GEN_21981); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22581 = 6'h11 == state ? $signed(digest_21) : $signed(_GEN_21982); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22582 = 6'h11 == state ? $signed(digest_22) : $signed(_GEN_21983); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22583 = 6'h11 == state ? $signed(digest_23) : $signed(_GEN_21984); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22584 = 6'h11 == state ? $signed(digest_24) : $signed(_GEN_21985); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22585 = 6'h11 == state ? $signed(digest_25) : $signed(_GEN_21986); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22586 = 6'h11 == state ? $signed(digest_26) : $signed(_GEN_21987); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22587 = 6'h11 == state ? $signed(digest_27) : $signed(_GEN_21988); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22588 = 6'h11 == state ? $signed(digest_28) : $signed(_GEN_21989); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22589 = 6'h11 == state ? $signed(digest_29) : $signed(_GEN_21990); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22590 = 6'h11 == state ? $signed(digest_30) : $signed(_GEN_21991); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22591 = 6'h11 == state ? $signed(digest_31) : $signed(_GEN_21992); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22592 = 6'h11 == state ? $signed(digest_32) : $signed(_GEN_21993); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22593 = 6'h11 == state ? $signed(digest_33) : $signed(_GEN_21994); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22594 = 6'h11 == state ? $signed(digest_34) : $signed(_GEN_21995); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22595 = 6'h11 == state ? $signed(digest_35) : $signed(_GEN_21996); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22596 = 6'h11 == state ? $signed(digest_36) : $signed(_GEN_21997); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22597 = 6'h11 == state ? $signed(digest_37) : $signed(_GEN_21998); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22598 = 6'h11 == state ? $signed(digest_38) : $signed(_GEN_21999); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22599 = 6'h11 == state ? $signed(digest_39) : $signed(_GEN_22000); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22600 = 6'h11 == state ? $signed(digest_40) : $signed(_GEN_22001); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22601 = 6'h11 == state ? $signed(digest_41) : $signed(_GEN_22002); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22602 = 6'h11 == state ? $signed(digest_42) : $signed(_GEN_22003); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22603 = 6'h11 == state ? $signed(digest_43) : $signed(_GEN_22004); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22604 = 6'h11 == state ? $signed(digest_44) : $signed(_GEN_22005); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22605 = 6'h11 == state ? $signed(digest_45) : $signed(_GEN_22006); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22606 = 6'h11 == state ? $signed(digest_46) : $signed(_GEN_22007); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22607 = 6'h11 == state ? $signed(digest_47) : $signed(_GEN_22008); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22608 = 6'h11 == state ? $signed(digest_48) : $signed(_GEN_22009); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22609 = 6'h11 == state ? $signed(digest_49) : $signed(_GEN_22010); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22610 = 6'h11 == state ? $signed(digest_50) : $signed(_GEN_22011); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22611 = 6'h11 == state ? $signed(digest_51) : $signed(_GEN_22012); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22612 = 6'h11 == state ? $signed(digest_52) : $signed(_GEN_22013); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22613 = 6'h11 == state ? $signed(digest_53) : $signed(_GEN_22014); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22614 = 6'h11 == state ? $signed(digest_54) : $signed(_GEN_22015); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22615 = 6'h11 == state ? $signed(digest_55) : $signed(_GEN_22016); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22616 = 6'h11 == state ? $signed(digest_56) : $signed(_GEN_22017); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22617 = 6'h11 == state ? $signed(digest_57) : $signed(_GEN_22018); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22618 = 6'h11 == state ? $signed(digest_58) : $signed(_GEN_22019); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22619 = 6'h11 == state ? $signed(digest_59) : $signed(_GEN_22020); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22620 = 6'h11 == state ? $signed(digest_60) : $signed(_GEN_22021); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22621 = 6'h11 == state ? $signed(digest_61) : $signed(_GEN_22022); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22622 = 6'h11 == state ? $signed(digest_62) : $signed(_GEN_22023); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22623 = 6'h11 == state ? $signed(digest_63) : $signed(_GEN_22024); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22624 = 6'h11 == state ? $signed(digest_64) : $signed(_GEN_22025); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22625 = 6'h11 == state ? $signed(digest_65) : $signed(_GEN_22026); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22626 = 6'h11 == state ? $signed(digest_66) : $signed(_GEN_22027); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22627 = 6'h11 == state ? $signed(digest_67) : $signed(_GEN_22028); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22628 = 6'h11 == state ? $signed(digest_68) : $signed(_GEN_22029); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22629 = 6'h11 == state ? $signed(digest_69) : $signed(_GEN_22030); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22630 = 6'h11 == state ? $signed(digest_70) : $signed(_GEN_22031); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22631 = 6'h11 == state ? $signed(digest_71) : $signed(_GEN_22032); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22632 = 6'h11 == state ? $signed(digest_72) : $signed(_GEN_22033); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22633 = 6'h11 == state ? $signed(digest_73) : $signed(_GEN_22034); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22634 = 6'h11 == state ? $signed(digest_74) : $signed(_GEN_22035); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22635 = 6'h11 == state ? $signed(digest_75) : $signed(_GEN_22036); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22636 = 6'h11 == state ? $signed(digest_76) : $signed(_GEN_22037); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22637 = 6'h11 == state ? $signed(digest_77) : $signed(_GEN_22038); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22638 = 6'h11 == state ? $signed(digest_78) : $signed(_GEN_22039); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_22639 = 6'h11 == state ? $signed(digest_79) : $signed(_GEN_22040); // @[digest.scala 81:19 53:21]
  wire  _GEN_22641 = 6'h11 == state ? 1'h0 : _GEN_22042; // @[digest.scala 81:19 58:25]
  wire  _GEN_22724 = 6'h11 == state ? 1'h0 : _GEN_22125; // @[digest.scala 81:19 63:25]
  wire  _GEN_22807 = 6'h11 == state ? 1'h0 : _GEN_22208; // @[digest.scala 81:19 68:25]
  wire  _GEN_22890 = 6'h11 == state ? 1'h0 : _GEN_22291; // @[digest.scala 81:19 73:25]
  wire  _GEN_22973 = 6'h11 == state ? 1'h0 : _GEN_22374; // @[digest.scala 81:19 78:25]
  wire [5:0] _GEN_22974 = 6'h10 == state ? _state_T_4 : _GEN_22376; // @[digest.scala 149:19 81:19]
  wire [31:0] _GEN_22975 = 6'h10 == state ? $signed(olda) : $signed(_GEN_22375); // @[digest.scala 29:19 81:19]
  wire [31:0] _GEN_22976 = 6'h10 == state ? $signed(oldb) : $signed(_GEN_22377); // @[digest.scala 30:19 81:19]
  wire [31:0] _GEN_22977 = 6'h10 == state ? $signed(oldc) : $signed(_GEN_22378); // @[digest.scala 31:19 81:19]
  wire [31:0] _GEN_22978 = 6'h10 == state ? $signed(oldd) : $signed(_GEN_22379); // @[digest.scala 32:19 81:19]
  wire [31:0] _GEN_22979 = 6'h10 == state ? $signed(olde) : $signed(_GEN_22380); // @[digest.scala 33:19 81:19]
  wire [31:0] _GEN_22980 = 6'h10 == state ? $signed(j) : $signed(_GEN_22381); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_22981 = 6'h10 == state ? $signed(w_0) : $signed(_GEN_22382); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22982 = 6'h10 == state ? $signed(w_1) : $signed(_GEN_22383); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22983 = 6'h10 == state ? $signed(w_2) : $signed(_GEN_22384); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22984 = 6'h10 == state ? $signed(w_3) : $signed(_GEN_22385); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22985 = 6'h10 == state ? $signed(w_4) : $signed(_GEN_22386); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22986 = 6'h10 == state ? $signed(w_5) : $signed(_GEN_22387); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22987 = 6'h10 == state ? $signed(w_6) : $signed(_GEN_22388); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22988 = 6'h10 == state ? $signed(w_7) : $signed(_GEN_22389); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22989 = 6'h10 == state ? $signed(w_8) : $signed(_GEN_22390); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22990 = 6'h10 == state ? $signed(w_9) : $signed(_GEN_22391); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22991 = 6'h10 == state ? $signed(w_10) : $signed(_GEN_22392); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22992 = 6'h10 == state ? $signed(w_11) : $signed(_GEN_22393); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22993 = 6'h10 == state ? $signed(w_12) : $signed(_GEN_22394); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22994 = 6'h10 == state ? $signed(w_13) : $signed(_GEN_22395); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22995 = 6'h10 == state ? $signed(w_14) : $signed(_GEN_22396); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22996 = 6'h10 == state ? $signed(w_15) : $signed(_GEN_22397); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22997 = 6'h10 == state ? $signed(w_16) : $signed(_GEN_22398); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22998 = 6'h10 == state ? $signed(w_17) : $signed(_GEN_22399); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_22999 = 6'h10 == state ? $signed(w_18) : $signed(_GEN_22400); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23000 = 6'h10 == state ? $signed(w_19) : $signed(_GEN_22401); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23001 = 6'h10 == state ? $signed(w_20) : $signed(_GEN_22402); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23002 = 6'h10 == state ? $signed(w_21) : $signed(_GEN_22403); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23003 = 6'h10 == state ? $signed(w_22) : $signed(_GEN_22404); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23004 = 6'h10 == state ? $signed(w_23) : $signed(_GEN_22405); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23005 = 6'h10 == state ? $signed(w_24) : $signed(_GEN_22406); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23006 = 6'h10 == state ? $signed(w_25) : $signed(_GEN_22407); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23007 = 6'h10 == state ? $signed(w_26) : $signed(_GEN_22408); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23008 = 6'h10 == state ? $signed(w_27) : $signed(_GEN_22409); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23009 = 6'h10 == state ? $signed(w_28) : $signed(_GEN_22410); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23010 = 6'h10 == state ? $signed(w_29) : $signed(_GEN_22411); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23011 = 6'h10 == state ? $signed(w_30) : $signed(_GEN_22412); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23012 = 6'h10 == state ? $signed(w_31) : $signed(_GEN_22413); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23013 = 6'h10 == state ? $signed(w_32) : $signed(_GEN_22414); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23014 = 6'h10 == state ? $signed(w_33) : $signed(_GEN_22415); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23015 = 6'h10 == state ? $signed(w_34) : $signed(_GEN_22416); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23016 = 6'h10 == state ? $signed(w_35) : $signed(_GEN_22417); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23017 = 6'h10 == state ? $signed(w_36) : $signed(_GEN_22418); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23018 = 6'h10 == state ? $signed(w_37) : $signed(_GEN_22419); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23019 = 6'h10 == state ? $signed(w_38) : $signed(_GEN_22420); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23020 = 6'h10 == state ? $signed(w_39) : $signed(_GEN_22421); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23021 = 6'h10 == state ? $signed(w_40) : $signed(_GEN_22422); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23022 = 6'h10 == state ? $signed(w_41) : $signed(_GEN_22423); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23023 = 6'h10 == state ? $signed(w_42) : $signed(_GEN_22424); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23024 = 6'h10 == state ? $signed(w_43) : $signed(_GEN_22425); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23025 = 6'h10 == state ? $signed(w_44) : $signed(_GEN_22426); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23026 = 6'h10 == state ? $signed(w_45) : $signed(_GEN_22427); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23027 = 6'h10 == state ? $signed(w_46) : $signed(_GEN_22428); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23028 = 6'h10 == state ? $signed(w_47) : $signed(_GEN_22429); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23029 = 6'h10 == state ? $signed(w_48) : $signed(_GEN_22430); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23030 = 6'h10 == state ? $signed(w_49) : $signed(_GEN_22431); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23031 = 6'h10 == state ? $signed(w_50) : $signed(_GEN_22432); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23032 = 6'h10 == state ? $signed(w_51) : $signed(_GEN_22433); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23033 = 6'h10 == state ? $signed(w_52) : $signed(_GEN_22434); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23034 = 6'h10 == state ? $signed(w_53) : $signed(_GEN_22435); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23035 = 6'h10 == state ? $signed(w_54) : $signed(_GEN_22436); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23036 = 6'h10 == state ? $signed(w_55) : $signed(_GEN_22437); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23037 = 6'h10 == state ? $signed(w_56) : $signed(_GEN_22438); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23038 = 6'h10 == state ? $signed(w_57) : $signed(_GEN_22439); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23039 = 6'h10 == state ? $signed(w_58) : $signed(_GEN_22440); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23040 = 6'h10 == state ? $signed(w_59) : $signed(_GEN_22441); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23041 = 6'h10 == state ? $signed(w_60) : $signed(_GEN_22442); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23042 = 6'h10 == state ? $signed(w_61) : $signed(_GEN_22443); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23043 = 6'h10 == state ? $signed(w_62) : $signed(_GEN_22444); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23044 = 6'h10 == state ? $signed(w_63) : $signed(_GEN_22445); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23045 = 6'h10 == state ? $signed(w_64) : $signed(_GEN_22446); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23046 = 6'h10 == state ? $signed(w_65) : $signed(_GEN_22447); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23047 = 6'h10 == state ? $signed(w_66) : $signed(_GEN_22448); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23048 = 6'h10 == state ? $signed(w_67) : $signed(_GEN_22449); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23049 = 6'h10 == state ? $signed(w_68) : $signed(_GEN_22450); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23050 = 6'h10 == state ? $signed(w_69) : $signed(_GEN_22451); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23051 = 6'h10 == state ? $signed(w_70) : $signed(_GEN_22452); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23052 = 6'h10 == state ? $signed(w_71) : $signed(_GEN_22453); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23053 = 6'h10 == state ? $signed(w_72) : $signed(_GEN_22454); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23054 = 6'h10 == state ? $signed(w_73) : $signed(_GEN_22455); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23055 = 6'h10 == state ? $signed(w_74) : $signed(_GEN_22456); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23056 = 6'h10 == state ? $signed(w_75) : $signed(_GEN_22457); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23057 = 6'h10 == state ? $signed(w_76) : $signed(_GEN_22458); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23058 = 6'h10 == state ? $signed(w_77) : $signed(_GEN_22459); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23059 = 6'h10 == state ? $signed(w_78) : $signed(_GEN_22460); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23060 = 6'h10 == state ? $signed(w_79) : $signed(_GEN_22461); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23061 = 6'h10 == state ? $signed(temp) : $signed(_GEN_22462); // @[digest.scala 38:19 81:19]
  wire  _GEN_23062 = 6'h10 == state ? 1'h0 : _GEN_22463; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_23065 = 6'h10 == state ? $signed(t) : $signed(_GEN_22466); // @[digest.scala 35:16 81:19]
  wire  _GEN_23066 = 6'h10 == state ? 1'h0 : _GEN_22467; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_23069 = 6'h10 == state ? $signed(e) : $signed(_GEN_22470); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_23070 = 6'h10 == state ? $signed(d) : $signed(_GEN_22471); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_23071 = 6'h10 == state ? $signed(c) : $signed(_GEN_22472); // @[digest.scala 26:16 81:19]
  wire  _GEN_23072 = 6'h10 == state ? 1'h0 : _GEN_22473; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_23075 = 6'h10 == state ? $signed(b) : $signed(_GEN_22476); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_23076 = 6'h10 == state ? $signed(a) : $signed(_GEN_22477); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_23077 = 6'h10 == state ? $signed(i) : $signed(_GEN_22478); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_23159 = 6'h10 == state ? $signed(digest_0) : $signed(_GEN_22560); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23160 = 6'h10 == state ? $signed(digest_1) : $signed(_GEN_22561); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23161 = 6'h10 == state ? $signed(digest_2) : $signed(_GEN_22562); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23162 = 6'h10 == state ? $signed(digest_3) : $signed(_GEN_22563); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23163 = 6'h10 == state ? $signed(digest_4) : $signed(_GEN_22564); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23164 = 6'h10 == state ? $signed(digest_5) : $signed(_GEN_22565); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23165 = 6'h10 == state ? $signed(digest_6) : $signed(_GEN_22566); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23166 = 6'h10 == state ? $signed(digest_7) : $signed(_GEN_22567); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23167 = 6'h10 == state ? $signed(digest_8) : $signed(_GEN_22568); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23168 = 6'h10 == state ? $signed(digest_9) : $signed(_GEN_22569); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23169 = 6'h10 == state ? $signed(digest_10) : $signed(_GEN_22570); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23170 = 6'h10 == state ? $signed(digest_11) : $signed(_GEN_22571); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23171 = 6'h10 == state ? $signed(digest_12) : $signed(_GEN_22572); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23172 = 6'h10 == state ? $signed(digest_13) : $signed(_GEN_22573); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23173 = 6'h10 == state ? $signed(digest_14) : $signed(_GEN_22574); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23174 = 6'h10 == state ? $signed(digest_15) : $signed(_GEN_22575); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23175 = 6'h10 == state ? $signed(digest_16) : $signed(_GEN_22576); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23176 = 6'h10 == state ? $signed(digest_17) : $signed(_GEN_22577); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23177 = 6'h10 == state ? $signed(digest_18) : $signed(_GEN_22578); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23178 = 6'h10 == state ? $signed(digest_19) : $signed(_GEN_22579); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23179 = 6'h10 == state ? $signed(digest_20) : $signed(_GEN_22580); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23180 = 6'h10 == state ? $signed(digest_21) : $signed(_GEN_22581); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23181 = 6'h10 == state ? $signed(digest_22) : $signed(_GEN_22582); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23182 = 6'h10 == state ? $signed(digest_23) : $signed(_GEN_22583); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23183 = 6'h10 == state ? $signed(digest_24) : $signed(_GEN_22584); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23184 = 6'h10 == state ? $signed(digest_25) : $signed(_GEN_22585); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23185 = 6'h10 == state ? $signed(digest_26) : $signed(_GEN_22586); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23186 = 6'h10 == state ? $signed(digest_27) : $signed(_GEN_22587); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23187 = 6'h10 == state ? $signed(digest_28) : $signed(_GEN_22588); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23188 = 6'h10 == state ? $signed(digest_29) : $signed(_GEN_22589); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23189 = 6'h10 == state ? $signed(digest_30) : $signed(_GEN_22590); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23190 = 6'h10 == state ? $signed(digest_31) : $signed(_GEN_22591); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23191 = 6'h10 == state ? $signed(digest_32) : $signed(_GEN_22592); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23192 = 6'h10 == state ? $signed(digest_33) : $signed(_GEN_22593); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23193 = 6'h10 == state ? $signed(digest_34) : $signed(_GEN_22594); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23194 = 6'h10 == state ? $signed(digest_35) : $signed(_GEN_22595); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23195 = 6'h10 == state ? $signed(digest_36) : $signed(_GEN_22596); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23196 = 6'h10 == state ? $signed(digest_37) : $signed(_GEN_22597); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23197 = 6'h10 == state ? $signed(digest_38) : $signed(_GEN_22598); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23198 = 6'h10 == state ? $signed(digest_39) : $signed(_GEN_22599); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23199 = 6'h10 == state ? $signed(digest_40) : $signed(_GEN_22600); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23200 = 6'h10 == state ? $signed(digest_41) : $signed(_GEN_22601); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23201 = 6'h10 == state ? $signed(digest_42) : $signed(_GEN_22602); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23202 = 6'h10 == state ? $signed(digest_43) : $signed(_GEN_22603); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23203 = 6'h10 == state ? $signed(digest_44) : $signed(_GEN_22604); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23204 = 6'h10 == state ? $signed(digest_45) : $signed(_GEN_22605); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23205 = 6'h10 == state ? $signed(digest_46) : $signed(_GEN_22606); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23206 = 6'h10 == state ? $signed(digest_47) : $signed(_GEN_22607); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23207 = 6'h10 == state ? $signed(digest_48) : $signed(_GEN_22608); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23208 = 6'h10 == state ? $signed(digest_49) : $signed(_GEN_22609); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23209 = 6'h10 == state ? $signed(digest_50) : $signed(_GEN_22610); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23210 = 6'h10 == state ? $signed(digest_51) : $signed(_GEN_22611); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23211 = 6'h10 == state ? $signed(digest_52) : $signed(_GEN_22612); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23212 = 6'h10 == state ? $signed(digest_53) : $signed(_GEN_22613); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23213 = 6'h10 == state ? $signed(digest_54) : $signed(_GEN_22614); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23214 = 6'h10 == state ? $signed(digest_55) : $signed(_GEN_22615); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23215 = 6'h10 == state ? $signed(digest_56) : $signed(_GEN_22616); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23216 = 6'h10 == state ? $signed(digest_57) : $signed(_GEN_22617); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23217 = 6'h10 == state ? $signed(digest_58) : $signed(_GEN_22618); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23218 = 6'h10 == state ? $signed(digest_59) : $signed(_GEN_22619); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23219 = 6'h10 == state ? $signed(digest_60) : $signed(_GEN_22620); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23220 = 6'h10 == state ? $signed(digest_61) : $signed(_GEN_22621); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23221 = 6'h10 == state ? $signed(digest_62) : $signed(_GEN_22622); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23222 = 6'h10 == state ? $signed(digest_63) : $signed(_GEN_22623); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23223 = 6'h10 == state ? $signed(digest_64) : $signed(_GEN_22624); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23224 = 6'h10 == state ? $signed(digest_65) : $signed(_GEN_22625); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23225 = 6'h10 == state ? $signed(digest_66) : $signed(_GEN_22626); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23226 = 6'h10 == state ? $signed(digest_67) : $signed(_GEN_22627); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23227 = 6'h10 == state ? $signed(digest_68) : $signed(_GEN_22628); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23228 = 6'h10 == state ? $signed(digest_69) : $signed(_GEN_22629); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23229 = 6'h10 == state ? $signed(digest_70) : $signed(_GEN_22630); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23230 = 6'h10 == state ? $signed(digest_71) : $signed(_GEN_22631); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23231 = 6'h10 == state ? $signed(digest_72) : $signed(_GEN_22632); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23232 = 6'h10 == state ? $signed(digest_73) : $signed(_GEN_22633); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23233 = 6'h10 == state ? $signed(digest_74) : $signed(_GEN_22634); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23234 = 6'h10 == state ? $signed(digest_75) : $signed(_GEN_22635); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23235 = 6'h10 == state ? $signed(digest_76) : $signed(_GEN_22636); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23236 = 6'h10 == state ? $signed(digest_77) : $signed(_GEN_22637); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23237 = 6'h10 == state ? $signed(digest_78) : $signed(_GEN_22638); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23238 = 6'h10 == state ? $signed(digest_79) : $signed(_GEN_22639); // @[digest.scala 81:19 53:21]
  wire  _GEN_23240 = 6'h10 == state ? 1'h0 : _GEN_22641; // @[digest.scala 81:19 58:25]
  wire  _GEN_23323 = 6'h10 == state ? 1'h0 : _GEN_22724; // @[digest.scala 81:19 63:25]
  wire  _GEN_23406 = 6'h10 == state ? 1'h0 : _GEN_22807; // @[digest.scala 81:19 68:25]
  wire  _GEN_23489 = 6'h10 == state ? 1'h0 : _GEN_22890; // @[digest.scala 81:19 73:25]
  wire  _GEN_23572 = 6'h10 == state ? 1'h0 : _GEN_22973; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_23573 = 6'hf == state ? $signed(32'sh0) : $signed(_GEN_23077); // @[digest.scala 145:15 81:19]
  wire [5:0] _GEN_23574 = 6'hf == state ? 6'h10 : _GEN_22974; // @[digest.scala 146:19 81:19]
  wire [31:0] _GEN_23575 = 6'hf == state ? $signed(olda) : $signed(_GEN_22975); // @[digest.scala 29:19 81:19]
  wire [31:0] _GEN_23576 = 6'hf == state ? $signed(oldb) : $signed(_GEN_22976); // @[digest.scala 30:19 81:19]
  wire [31:0] _GEN_23577 = 6'hf == state ? $signed(oldc) : $signed(_GEN_22977); // @[digest.scala 31:19 81:19]
  wire [31:0] _GEN_23578 = 6'hf == state ? $signed(oldd) : $signed(_GEN_22978); // @[digest.scala 32:19 81:19]
  wire [31:0] _GEN_23579 = 6'hf == state ? $signed(olde) : $signed(_GEN_22979); // @[digest.scala 33:19 81:19]
  wire [31:0] _GEN_23580 = 6'hf == state ? $signed(j) : $signed(_GEN_22980); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_23581 = 6'hf == state ? $signed(w_0) : $signed(_GEN_22981); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23582 = 6'hf == state ? $signed(w_1) : $signed(_GEN_22982); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23583 = 6'hf == state ? $signed(w_2) : $signed(_GEN_22983); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23584 = 6'hf == state ? $signed(w_3) : $signed(_GEN_22984); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23585 = 6'hf == state ? $signed(w_4) : $signed(_GEN_22985); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23586 = 6'hf == state ? $signed(w_5) : $signed(_GEN_22986); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23587 = 6'hf == state ? $signed(w_6) : $signed(_GEN_22987); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23588 = 6'hf == state ? $signed(w_7) : $signed(_GEN_22988); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23589 = 6'hf == state ? $signed(w_8) : $signed(_GEN_22989); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23590 = 6'hf == state ? $signed(w_9) : $signed(_GEN_22990); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23591 = 6'hf == state ? $signed(w_10) : $signed(_GEN_22991); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23592 = 6'hf == state ? $signed(w_11) : $signed(_GEN_22992); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23593 = 6'hf == state ? $signed(w_12) : $signed(_GEN_22993); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23594 = 6'hf == state ? $signed(w_13) : $signed(_GEN_22994); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23595 = 6'hf == state ? $signed(w_14) : $signed(_GEN_22995); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23596 = 6'hf == state ? $signed(w_15) : $signed(_GEN_22996); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23597 = 6'hf == state ? $signed(w_16) : $signed(_GEN_22997); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23598 = 6'hf == state ? $signed(w_17) : $signed(_GEN_22998); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23599 = 6'hf == state ? $signed(w_18) : $signed(_GEN_22999); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23600 = 6'hf == state ? $signed(w_19) : $signed(_GEN_23000); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23601 = 6'hf == state ? $signed(w_20) : $signed(_GEN_23001); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23602 = 6'hf == state ? $signed(w_21) : $signed(_GEN_23002); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23603 = 6'hf == state ? $signed(w_22) : $signed(_GEN_23003); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23604 = 6'hf == state ? $signed(w_23) : $signed(_GEN_23004); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23605 = 6'hf == state ? $signed(w_24) : $signed(_GEN_23005); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23606 = 6'hf == state ? $signed(w_25) : $signed(_GEN_23006); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23607 = 6'hf == state ? $signed(w_26) : $signed(_GEN_23007); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23608 = 6'hf == state ? $signed(w_27) : $signed(_GEN_23008); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23609 = 6'hf == state ? $signed(w_28) : $signed(_GEN_23009); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23610 = 6'hf == state ? $signed(w_29) : $signed(_GEN_23010); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23611 = 6'hf == state ? $signed(w_30) : $signed(_GEN_23011); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23612 = 6'hf == state ? $signed(w_31) : $signed(_GEN_23012); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23613 = 6'hf == state ? $signed(w_32) : $signed(_GEN_23013); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23614 = 6'hf == state ? $signed(w_33) : $signed(_GEN_23014); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23615 = 6'hf == state ? $signed(w_34) : $signed(_GEN_23015); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23616 = 6'hf == state ? $signed(w_35) : $signed(_GEN_23016); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23617 = 6'hf == state ? $signed(w_36) : $signed(_GEN_23017); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23618 = 6'hf == state ? $signed(w_37) : $signed(_GEN_23018); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23619 = 6'hf == state ? $signed(w_38) : $signed(_GEN_23019); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23620 = 6'hf == state ? $signed(w_39) : $signed(_GEN_23020); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23621 = 6'hf == state ? $signed(w_40) : $signed(_GEN_23021); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23622 = 6'hf == state ? $signed(w_41) : $signed(_GEN_23022); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23623 = 6'hf == state ? $signed(w_42) : $signed(_GEN_23023); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23624 = 6'hf == state ? $signed(w_43) : $signed(_GEN_23024); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23625 = 6'hf == state ? $signed(w_44) : $signed(_GEN_23025); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23626 = 6'hf == state ? $signed(w_45) : $signed(_GEN_23026); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23627 = 6'hf == state ? $signed(w_46) : $signed(_GEN_23027); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23628 = 6'hf == state ? $signed(w_47) : $signed(_GEN_23028); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23629 = 6'hf == state ? $signed(w_48) : $signed(_GEN_23029); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23630 = 6'hf == state ? $signed(w_49) : $signed(_GEN_23030); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23631 = 6'hf == state ? $signed(w_50) : $signed(_GEN_23031); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23632 = 6'hf == state ? $signed(w_51) : $signed(_GEN_23032); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23633 = 6'hf == state ? $signed(w_52) : $signed(_GEN_23033); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23634 = 6'hf == state ? $signed(w_53) : $signed(_GEN_23034); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23635 = 6'hf == state ? $signed(w_54) : $signed(_GEN_23035); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23636 = 6'hf == state ? $signed(w_55) : $signed(_GEN_23036); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23637 = 6'hf == state ? $signed(w_56) : $signed(_GEN_23037); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23638 = 6'hf == state ? $signed(w_57) : $signed(_GEN_23038); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23639 = 6'hf == state ? $signed(w_58) : $signed(_GEN_23039); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23640 = 6'hf == state ? $signed(w_59) : $signed(_GEN_23040); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23641 = 6'hf == state ? $signed(w_60) : $signed(_GEN_23041); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23642 = 6'hf == state ? $signed(w_61) : $signed(_GEN_23042); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23643 = 6'hf == state ? $signed(w_62) : $signed(_GEN_23043); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23644 = 6'hf == state ? $signed(w_63) : $signed(_GEN_23044); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23645 = 6'hf == state ? $signed(w_64) : $signed(_GEN_23045); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23646 = 6'hf == state ? $signed(w_65) : $signed(_GEN_23046); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23647 = 6'hf == state ? $signed(w_66) : $signed(_GEN_23047); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23648 = 6'hf == state ? $signed(w_67) : $signed(_GEN_23048); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23649 = 6'hf == state ? $signed(w_68) : $signed(_GEN_23049); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23650 = 6'hf == state ? $signed(w_69) : $signed(_GEN_23050); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23651 = 6'hf == state ? $signed(w_70) : $signed(_GEN_23051); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23652 = 6'hf == state ? $signed(w_71) : $signed(_GEN_23052); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23653 = 6'hf == state ? $signed(w_72) : $signed(_GEN_23053); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23654 = 6'hf == state ? $signed(w_73) : $signed(_GEN_23054); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23655 = 6'hf == state ? $signed(w_74) : $signed(_GEN_23055); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23656 = 6'hf == state ? $signed(w_75) : $signed(_GEN_23056); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23657 = 6'hf == state ? $signed(w_76) : $signed(_GEN_23057); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23658 = 6'hf == state ? $signed(w_77) : $signed(_GEN_23058); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23659 = 6'hf == state ? $signed(w_78) : $signed(_GEN_23059); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23660 = 6'hf == state ? $signed(w_79) : $signed(_GEN_23060); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_23661 = 6'hf == state ? $signed(temp) : $signed(_GEN_23061); // @[digest.scala 38:19 81:19]
  wire  _GEN_23662 = 6'hf == state ? 1'h0 : _GEN_23062; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_23665 = 6'hf == state ? $signed(t) : $signed(_GEN_23065); // @[digest.scala 35:16 81:19]
  wire  _GEN_23666 = 6'hf == state ? 1'h0 : _GEN_23066; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_23669 = 6'hf == state ? $signed(e) : $signed(_GEN_23069); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_23670 = 6'hf == state ? $signed(d) : $signed(_GEN_23070); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_23671 = 6'hf == state ? $signed(c) : $signed(_GEN_23071); // @[digest.scala 26:16 81:19]
  wire  _GEN_23672 = 6'hf == state ? 1'h0 : _GEN_23072; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_23675 = 6'hf == state ? $signed(b) : $signed(_GEN_23075); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_23676 = 6'hf == state ? $signed(a) : $signed(_GEN_23076); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_23758 = 6'hf == state ? $signed(digest_0) : $signed(_GEN_23159); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23759 = 6'hf == state ? $signed(digest_1) : $signed(_GEN_23160); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23760 = 6'hf == state ? $signed(digest_2) : $signed(_GEN_23161); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23761 = 6'hf == state ? $signed(digest_3) : $signed(_GEN_23162); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23762 = 6'hf == state ? $signed(digest_4) : $signed(_GEN_23163); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23763 = 6'hf == state ? $signed(digest_5) : $signed(_GEN_23164); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23764 = 6'hf == state ? $signed(digest_6) : $signed(_GEN_23165); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23765 = 6'hf == state ? $signed(digest_7) : $signed(_GEN_23166); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23766 = 6'hf == state ? $signed(digest_8) : $signed(_GEN_23167); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23767 = 6'hf == state ? $signed(digest_9) : $signed(_GEN_23168); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23768 = 6'hf == state ? $signed(digest_10) : $signed(_GEN_23169); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23769 = 6'hf == state ? $signed(digest_11) : $signed(_GEN_23170); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23770 = 6'hf == state ? $signed(digest_12) : $signed(_GEN_23171); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23771 = 6'hf == state ? $signed(digest_13) : $signed(_GEN_23172); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23772 = 6'hf == state ? $signed(digest_14) : $signed(_GEN_23173); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23773 = 6'hf == state ? $signed(digest_15) : $signed(_GEN_23174); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23774 = 6'hf == state ? $signed(digest_16) : $signed(_GEN_23175); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23775 = 6'hf == state ? $signed(digest_17) : $signed(_GEN_23176); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23776 = 6'hf == state ? $signed(digest_18) : $signed(_GEN_23177); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23777 = 6'hf == state ? $signed(digest_19) : $signed(_GEN_23178); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23778 = 6'hf == state ? $signed(digest_20) : $signed(_GEN_23179); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23779 = 6'hf == state ? $signed(digest_21) : $signed(_GEN_23180); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23780 = 6'hf == state ? $signed(digest_22) : $signed(_GEN_23181); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23781 = 6'hf == state ? $signed(digest_23) : $signed(_GEN_23182); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23782 = 6'hf == state ? $signed(digest_24) : $signed(_GEN_23183); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23783 = 6'hf == state ? $signed(digest_25) : $signed(_GEN_23184); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23784 = 6'hf == state ? $signed(digest_26) : $signed(_GEN_23185); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23785 = 6'hf == state ? $signed(digest_27) : $signed(_GEN_23186); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23786 = 6'hf == state ? $signed(digest_28) : $signed(_GEN_23187); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23787 = 6'hf == state ? $signed(digest_29) : $signed(_GEN_23188); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23788 = 6'hf == state ? $signed(digest_30) : $signed(_GEN_23189); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23789 = 6'hf == state ? $signed(digest_31) : $signed(_GEN_23190); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23790 = 6'hf == state ? $signed(digest_32) : $signed(_GEN_23191); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23791 = 6'hf == state ? $signed(digest_33) : $signed(_GEN_23192); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23792 = 6'hf == state ? $signed(digest_34) : $signed(_GEN_23193); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23793 = 6'hf == state ? $signed(digest_35) : $signed(_GEN_23194); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23794 = 6'hf == state ? $signed(digest_36) : $signed(_GEN_23195); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23795 = 6'hf == state ? $signed(digest_37) : $signed(_GEN_23196); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23796 = 6'hf == state ? $signed(digest_38) : $signed(_GEN_23197); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23797 = 6'hf == state ? $signed(digest_39) : $signed(_GEN_23198); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23798 = 6'hf == state ? $signed(digest_40) : $signed(_GEN_23199); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23799 = 6'hf == state ? $signed(digest_41) : $signed(_GEN_23200); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23800 = 6'hf == state ? $signed(digest_42) : $signed(_GEN_23201); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23801 = 6'hf == state ? $signed(digest_43) : $signed(_GEN_23202); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23802 = 6'hf == state ? $signed(digest_44) : $signed(_GEN_23203); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23803 = 6'hf == state ? $signed(digest_45) : $signed(_GEN_23204); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23804 = 6'hf == state ? $signed(digest_46) : $signed(_GEN_23205); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23805 = 6'hf == state ? $signed(digest_47) : $signed(_GEN_23206); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23806 = 6'hf == state ? $signed(digest_48) : $signed(_GEN_23207); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23807 = 6'hf == state ? $signed(digest_49) : $signed(_GEN_23208); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23808 = 6'hf == state ? $signed(digest_50) : $signed(_GEN_23209); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23809 = 6'hf == state ? $signed(digest_51) : $signed(_GEN_23210); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23810 = 6'hf == state ? $signed(digest_52) : $signed(_GEN_23211); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23811 = 6'hf == state ? $signed(digest_53) : $signed(_GEN_23212); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23812 = 6'hf == state ? $signed(digest_54) : $signed(_GEN_23213); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23813 = 6'hf == state ? $signed(digest_55) : $signed(_GEN_23214); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23814 = 6'hf == state ? $signed(digest_56) : $signed(_GEN_23215); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23815 = 6'hf == state ? $signed(digest_57) : $signed(_GEN_23216); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23816 = 6'hf == state ? $signed(digest_58) : $signed(_GEN_23217); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23817 = 6'hf == state ? $signed(digest_59) : $signed(_GEN_23218); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23818 = 6'hf == state ? $signed(digest_60) : $signed(_GEN_23219); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23819 = 6'hf == state ? $signed(digest_61) : $signed(_GEN_23220); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23820 = 6'hf == state ? $signed(digest_62) : $signed(_GEN_23221); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23821 = 6'hf == state ? $signed(digest_63) : $signed(_GEN_23222); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23822 = 6'hf == state ? $signed(digest_64) : $signed(_GEN_23223); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23823 = 6'hf == state ? $signed(digest_65) : $signed(_GEN_23224); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23824 = 6'hf == state ? $signed(digest_66) : $signed(_GEN_23225); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23825 = 6'hf == state ? $signed(digest_67) : $signed(_GEN_23226); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23826 = 6'hf == state ? $signed(digest_68) : $signed(_GEN_23227); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23827 = 6'hf == state ? $signed(digest_69) : $signed(_GEN_23228); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23828 = 6'hf == state ? $signed(digest_70) : $signed(_GEN_23229); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23829 = 6'hf == state ? $signed(digest_71) : $signed(_GEN_23230); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23830 = 6'hf == state ? $signed(digest_72) : $signed(_GEN_23231); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23831 = 6'hf == state ? $signed(digest_73) : $signed(_GEN_23232); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23832 = 6'hf == state ? $signed(digest_74) : $signed(_GEN_23233); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23833 = 6'hf == state ? $signed(digest_75) : $signed(_GEN_23234); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23834 = 6'hf == state ? $signed(digest_76) : $signed(_GEN_23235); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23835 = 6'hf == state ? $signed(digest_77) : $signed(_GEN_23236); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23836 = 6'hf == state ? $signed(digest_78) : $signed(_GEN_23237); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_23837 = 6'hf == state ? $signed(digest_79) : $signed(_GEN_23238); // @[digest.scala 81:19 53:21]
  wire  _GEN_23839 = 6'hf == state ? 1'h0 : _GEN_23240; // @[digest.scala 81:19 58:25]
  wire  _GEN_23922 = 6'hf == state ? 1'h0 : _GEN_23323; // @[digest.scala 81:19 63:25]
  wire  _GEN_24005 = 6'hf == state ? 1'h0 : _GEN_23406; // @[digest.scala 81:19 68:25]
  wire  _GEN_24088 = 6'hf == state ? 1'h0 : _GEN_23489; // @[digest.scala 81:19 73:25]
  wire  _GEN_24171 = 6'hf == state ? 1'h0 : _GEN_23572; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_24172 = 6'he == state ? $signed(-32'sh3c2d1e10) : $signed(_GEN_23669); // @[digest.scala 141:15 81:19]
  wire [5:0] _GEN_24173 = 6'he == state ? 6'hf : _GEN_23574; // @[digest.scala 142:19 81:19]
  wire [31:0] _GEN_24174 = 6'he == state ? $signed(i) : $signed(_GEN_23573); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_24175 = 6'he == state ? $signed(olda) : $signed(_GEN_23575); // @[digest.scala 29:19 81:19]
  wire [31:0] _GEN_24176 = 6'he == state ? $signed(oldb) : $signed(_GEN_23576); // @[digest.scala 30:19 81:19]
  wire [31:0] _GEN_24177 = 6'he == state ? $signed(oldc) : $signed(_GEN_23577); // @[digest.scala 31:19 81:19]
  wire [31:0] _GEN_24178 = 6'he == state ? $signed(oldd) : $signed(_GEN_23578); // @[digest.scala 32:19 81:19]
  wire [31:0] _GEN_24179 = 6'he == state ? $signed(olde) : $signed(_GEN_23579); // @[digest.scala 33:19 81:19]
  wire [31:0] _GEN_24180 = 6'he == state ? $signed(j) : $signed(_GEN_23580); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_24181 = 6'he == state ? $signed(w_0) : $signed(_GEN_23581); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24182 = 6'he == state ? $signed(w_1) : $signed(_GEN_23582); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24183 = 6'he == state ? $signed(w_2) : $signed(_GEN_23583); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24184 = 6'he == state ? $signed(w_3) : $signed(_GEN_23584); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24185 = 6'he == state ? $signed(w_4) : $signed(_GEN_23585); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24186 = 6'he == state ? $signed(w_5) : $signed(_GEN_23586); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24187 = 6'he == state ? $signed(w_6) : $signed(_GEN_23587); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24188 = 6'he == state ? $signed(w_7) : $signed(_GEN_23588); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24189 = 6'he == state ? $signed(w_8) : $signed(_GEN_23589); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24190 = 6'he == state ? $signed(w_9) : $signed(_GEN_23590); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24191 = 6'he == state ? $signed(w_10) : $signed(_GEN_23591); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24192 = 6'he == state ? $signed(w_11) : $signed(_GEN_23592); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24193 = 6'he == state ? $signed(w_12) : $signed(_GEN_23593); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24194 = 6'he == state ? $signed(w_13) : $signed(_GEN_23594); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24195 = 6'he == state ? $signed(w_14) : $signed(_GEN_23595); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24196 = 6'he == state ? $signed(w_15) : $signed(_GEN_23596); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24197 = 6'he == state ? $signed(w_16) : $signed(_GEN_23597); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24198 = 6'he == state ? $signed(w_17) : $signed(_GEN_23598); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24199 = 6'he == state ? $signed(w_18) : $signed(_GEN_23599); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24200 = 6'he == state ? $signed(w_19) : $signed(_GEN_23600); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24201 = 6'he == state ? $signed(w_20) : $signed(_GEN_23601); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24202 = 6'he == state ? $signed(w_21) : $signed(_GEN_23602); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24203 = 6'he == state ? $signed(w_22) : $signed(_GEN_23603); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24204 = 6'he == state ? $signed(w_23) : $signed(_GEN_23604); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24205 = 6'he == state ? $signed(w_24) : $signed(_GEN_23605); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24206 = 6'he == state ? $signed(w_25) : $signed(_GEN_23606); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24207 = 6'he == state ? $signed(w_26) : $signed(_GEN_23607); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24208 = 6'he == state ? $signed(w_27) : $signed(_GEN_23608); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24209 = 6'he == state ? $signed(w_28) : $signed(_GEN_23609); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24210 = 6'he == state ? $signed(w_29) : $signed(_GEN_23610); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24211 = 6'he == state ? $signed(w_30) : $signed(_GEN_23611); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24212 = 6'he == state ? $signed(w_31) : $signed(_GEN_23612); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24213 = 6'he == state ? $signed(w_32) : $signed(_GEN_23613); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24214 = 6'he == state ? $signed(w_33) : $signed(_GEN_23614); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24215 = 6'he == state ? $signed(w_34) : $signed(_GEN_23615); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24216 = 6'he == state ? $signed(w_35) : $signed(_GEN_23616); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24217 = 6'he == state ? $signed(w_36) : $signed(_GEN_23617); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24218 = 6'he == state ? $signed(w_37) : $signed(_GEN_23618); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24219 = 6'he == state ? $signed(w_38) : $signed(_GEN_23619); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24220 = 6'he == state ? $signed(w_39) : $signed(_GEN_23620); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24221 = 6'he == state ? $signed(w_40) : $signed(_GEN_23621); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24222 = 6'he == state ? $signed(w_41) : $signed(_GEN_23622); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24223 = 6'he == state ? $signed(w_42) : $signed(_GEN_23623); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24224 = 6'he == state ? $signed(w_43) : $signed(_GEN_23624); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24225 = 6'he == state ? $signed(w_44) : $signed(_GEN_23625); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24226 = 6'he == state ? $signed(w_45) : $signed(_GEN_23626); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24227 = 6'he == state ? $signed(w_46) : $signed(_GEN_23627); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24228 = 6'he == state ? $signed(w_47) : $signed(_GEN_23628); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24229 = 6'he == state ? $signed(w_48) : $signed(_GEN_23629); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24230 = 6'he == state ? $signed(w_49) : $signed(_GEN_23630); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24231 = 6'he == state ? $signed(w_50) : $signed(_GEN_23631); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24232 = 6'he == state ? $signed(w_51) : $signed(_GEN_23632); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24233 = 6'he == state ? $signed(w_52) : $signed(_GEN_23633); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24234 = 6'he == state ? $signed(w_53) : $signed(_GEN_23634); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24235 = 6'he == state ? $signed(w_54) : $signed(_GEN_23635); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24236 = 6'he == state ? $signed(w_55) : $signed(_GEN_23636); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24237 = 6'he == state ? $signed(w_56) : $signed(_GEN_23637); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24238 = 6'he == state ? $signed(w_57) : $signed(_GEN_23638); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24239 = 6'he == state ? $signed(w_58) : $signed(_GEN_23639); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24240 = 6'he == state ? $signed(w_59) : $signed(_GEN_23640); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24241 = 6'he == state ? $signed(w_60) : $signed(_GEN_23641); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24242 = 6'he == state ? $signed(w_61) : $signed(_GEN_23642); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24243 = 6'he == state ? $signed(w_62) : $signed(_GEN_23643); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24244 = 6'he == state ? $signed(w_63) : $signed(_GEN_23644); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24245 = 6'he == state ? $signed(w_64) : $signed(_GEN_23645); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24246 = 6'he == state ? $signed(w_65) : $signed(_GEN_23646); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24247 = 6'he == state ? $signed(w_66) : $signed(_GEN_23647); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24248 = 6'he == state ? $signed(w_67) : $signed(_GEN_23648); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24249 = 6'he == state ? $signed(w_68) : $signed(_GEN_23649); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24250 = 6'he == state ? $signed(w_69) : $signed(_GEN_23650); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24251 = 6'he == state ? $signed(w_70) : $signed(_GEN_23651); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24252 = 6'he == state ? $signed(w_71) : $signed(_GEN_23652); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24253 = 6'he == state ? $signed(w_72) : $signed(_GEN_23653); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24254 = 6'he == state ? $signed(w_73) : $signed(_GEN_23654); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24255 = 6'he == state ? $signed(w_74) : $signed(_GEN_23655); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24256 = 6'he == state ? $signed(w_75) : $signed(_GEN_23656); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24257 = 6'he == state ? $signed(w_76) : $signed(_GEN_23657); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24258 = 6'he == state ? $signed(w_77) : $signed(_GEN_23658); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24259 = 6'he == state ? $signed(w_78) : $signed(_GEN_23659); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24260 = 6'he == state ? $signed(w_79) : $signed(_GEN_23660); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24261 = 6'he == state ? $signed(temp) : $signed(_GEN_23661); // @[digest.scala 38:19 81:19]
  wire  _GEN_24262 = 6'he == state ? 1'h0 : _GEN_23662; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_24265 = 6'he == state ? $signed(t) : $signed(_GEN_23665); // @[digest.scala 35:16 81:19]
  wire  _GEN_24266 = 6'he == state ? 1'h0 : _GEN_23666; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_24269 = 6'he == state ? $signed(d) : $signed(_GEN_23670); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_24270 = 6'he == state ? $signed(c) : $signed(_GEN_23671); // @[digest.scala 26:16 81:19]
  wire  _GEN_24271 = 6'he == state ? 1'h0 : _GEN_23672; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_24274 = 6'he == state ? $signed(b) : $signed(_GEN_23675); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_24275 = 6'he == state ? $signed(a) : $signed(_GEN_23676); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_24357 = 6'he == state ? $signed(digest_0) : $signed(_GEN_23758); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24358 = 6'he == state ? $signed(digest_1) : $signed(_GEN_23759); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24359 = 6'he == state ? $signed(digest_2) : $signed(_GEN_23760); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24360 = 6'he == state ? $signed(digest_3) : $signed(_GEN_23761); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24361 = 6'he == state ? $signed(digest_4) : $signed(_GEN_23762); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24362 = 6'he == state ? $signed(digest_5) : $signed(_GEN_23763); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24363 = 6'he == state ? $signed(digest_6) : $signed(_GEN_23764); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24364 = 6'he == state ? $signed(digest_7) : $signed(_GEN_23765); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24365 = 6'he == state ? $signed(digest_8) : $signed(_GEN_23766); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24366 = 6'he == state ? $signed(digest_9) : $signed(_GEN_23767); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24367 = 6'he == state ? $signed(digest_10) : $signed(_GEN_23768); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24368 = 6'he == state ? $signed(digest_11) : $signed(_GEN_23769); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24369 = 6'he == state ? $signed(digest_12) : $signed(_GEN_23770); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24370 = 6'he == state ? $signed(digest_13) : $signed(_GEN_23771); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24371 = 6'he == state ? $signed(digest_14) : $signed(_GEN_23772); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24372 = 6'he == state ? $signed(digest_15) : $signed(_GEN_23773); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24373 = 6'he == state ? $signed(digest_16) : $signed(_GEN_23774); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24374 = 6'he == state ? $signed(digest_17) : $signed(_GEN_23775); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24375 = 6'he == state ? $signed(digest_18) : $signed(_GEN_23776); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24376 = 6'he == state ? $signed(digest_19) : $signed(_GEN_23777); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24377 = 6'he == state ? $signed(digest_20) : $signed(_GEN_23778); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24378 = 6'he == state ? $signed(digest_21) : $signed(_GEN_23779); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24379 = 6'he == state ? $signed(digest_22) : $signed(_GEN_23780); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24380 = 6'he == state ? $signed(digest_23) : $signed(_GEN_23781); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24381 = 6'he == state ? $signed(digest_24) : $signed(_GEN_23782); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24382 = 6'he == state ? $signed(digest_25) : $signed(_GEN_23783); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24383 = 6'he == state ? $signed(digest_26) : $signed(_GEN_23784); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24384 = 6'he == state ? $signed(digest_27) : $signed(_GEN_23785); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24385 = 6'he == state ? $signed(digest_28) : $signed(_GEN_23786); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24386 = 6'he == state ? $signed(digest_29) : $signed(_GEN_23787); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24387 = 6'he == state ? $signed(digest_30) : $signed(_GEN_23788); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24388 = 6'he == state ? $signed(digest_31) : $signed(_GEN_23789); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24389 = 6'he == state ? $signed(digest_32) : $signed(_GEN_23790); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24390 = 6'he == state ? $signed(digest_33) : $signed(_GEN_23791); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24391 = 6'he == state ? $signed(digest_34) : $signed(_GEN_23792); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24392 = 6'he == state ? $signed(digest_35) : $signed(_GEN_23793); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24393 = 6'he == state ? $signed(digest_36) : $signed(_GEN_23794); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24394 = 6'he == state ? $signed(digest_37) : $signed(_GEN_23795); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24395 = 6'he == state ? $signed(digest_38) : $signed(_GEN_23796); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24396 = 6'he == state ? $signed(digest_39) : $signed(_GEN_23797); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24397 = 6'he == state ? $signed(digest_40) : $signed(_GEN_23798); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24398 = 6'he == state ? $signed(digest_41) : $signed(_GEN_23799); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24399 = 6'he == state ? $signed(digest_42) : $signed(_GEN_23800); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24400 = 6'he == state ? $signed(digest_43) : $signed(_GEN_23801); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24401 = 6'he == state ? $signed(digest_44) : $signed(_GEN_23802); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24402 = 6'he == state ? $signed(digest_45) : $signed(_GEN_23803); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24403 = 6'he == state ? $signed(digest_46) : $signed(_GEN_23804); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24404 = 6'he == state ? $signed(digest_47) : $signed(_GEN_23805); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24405 = 6'he == state ? $signed(digest_48) : $signed(_GEN_23806); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24406 = 6'he == state ? $signed(digest_49) : $signed(_GEN_23807); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24407 = 6'he == state ? $signed(digest_50) : $signed(_GEN_23808); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24408 = 6'he == state ? $signed(digest_51) : $signed(_GEN_23809); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24409 = 6'he == state ? $signed(digest_52) : $signed(_GEN_23810); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24410 = 6'he == state ? $signed(digest_53) : $signed(_GEN_23811); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24411 = 6'he == state ? $signed(digest_54) : $signed(_GEN_23812); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24412 = 6'he == state ? $signed(digest_55) : $signed(_GEN_23813); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24413 = 6'he == state ? $signed(digest_56) : $signed(_GEN_23814); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24414 = 6'he == state ? $signed(digest_57) : $signed(_GEN_23815); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24415 = 6'he == state ? $signed(digest_58) : $signed(_GEN_23816); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24416 = 6'he == state ? $signed(digest_59) : $signed(_GEN_23817); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24417 = 6'he == state ? $signed(digest_60) : $signed(_GEN_23818); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24418 = 6'he == state ? $signed(digest_61) : $signed(_GEN_23819); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24419 = 6'he == state ? $signed(digest_62) : $signed(_GEN_23820); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24420 = 6'he == state ? $signed(digest_63) : $signed(_GEN_23821); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24421 = 6'he == state ? $signed(digest_64) : $signed(_GEN_23822); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24422 = 6'he == state ? $signed(digest_65) : $signed(_GEN_23823); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24423 = 6'he == state ? $signed(digest_66) : $signed(_GEN_23824); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24424 = 6'he == state ? $signed(digest_67) : $signed(_GEN_23825); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24425 = 6'he == state ? $signed(digest_68) : $signed(_GEN_23826); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24426 = 6'he == state ? $signed(digest_69) : $signed(_GEN_23827); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24427 = 6'he == state ? $signed(digest_70) : $signed(_GEN_23828); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24428 = 6'he == state ? $signed(digest_71) : $signed(_GEN_23829); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24429 = 6'he == state ? $signed(digest_72) : $signed(_GEN_23830); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24430 = 6'he == state ? $signed(digest_73) : $signed(_GEN_23831); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24431 = 6'he == state ? $signed(digest_74) : $signed(_GEN_23832); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24432 = 6'he == state ? $signed(digest_75) : $signed(_GEN_23833); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24433 = 6'he == state ? $signed(digest_76) : $signed(_GEN_23834); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24434 = 6'he == state ? $signed(digest_77) : $signed(_GEN_23835); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24435 = 6'he == state ? $signed(digest_78) : $signed(_GEN_23836); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24436 = 6'he == state ? $signed(digest_79) : $signed(_GEN_23837); // @[digest.scala 81:19 53:21]
  wire  _GEN_24438 = 6'he == state ? 1'h0 : _GEN_23839; // @[digest.scala 81:19 58:25]
  wire  _GEN_24521 = 6'he == state ? 1'h0 : _GEN_23922; // @[digest.scala 81:19 63:25]
  wire  _GEN_24604 = 6'he == state ? 1'h0 : _GEN_24005; // @[digest.scala 81:19 68:25]
  wire  _GEN_24687 = 6'he == state ? 1'h0 : _GEN_24088; // @[digest.scala 81:19 73:25]
  wire  _GEN_24770 = 6'he == state ? 1'h0 : _GEN_24171; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_24771 = 6'hd == state ? $signed(32'sh10325476) : $signed(_GEN_24269); // @[digest.scala 137:15 81:19]
  wire [5:0] _GEN_24772 = 6'hd == state ? 6'he : _GEN_24173; // @[digest.scala 138:19 81:19]
  wire [31:0] _GEN_24773 = 6'hd == state ? $signed(e) : $signed(_GEN_24172); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_24774 = 6'hd == state ? $signed(i) : $signed(_GEN_24174); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_24775 = 6'hd == state ? $signed(olda) : $signed(_GEN_24175); // @[digest.scala 29:19 81:19]
  wire [31:0] _GEN_24776 = 6'hd == state ? $signed(oldb) : $signed(_GEN_24176); // @[digest.scala 30:19 81:19]
  wire [31:0] _GEN_24777 = 6'hd == state ? $signed(oldc) : $signed(_GEN_24177); // @[digest.scala 31:19 81:19]
  wire [31:0] _GEN_24778 = 6'hd == state ? $signed(oldd) : $signed(_GEN_24178); // @[digest.scala 32:19 81:19]
  wire [31:0] _GEN_24779 = 6'hd == state ? $signed(olde) : $signed(_GEN_24179); // @[digest.scala 33:19 81:19]
  wire [31:0] _GEN_24780 = 6'hd == state ? $signed(j) : $signed(_GEN_24180); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_24781 = 6'hd == state ? $signed(w_0) : $signed(_GEN_24181); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24782 = 6'hd == state ? $signed(w_1) : $signed(_GEN_24182); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24783 = 6'hd == state ? $signed(w_2) : $signed(_GEN_24183); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24784 = 6'hd == state ? $signed(w_3) : $signed(_GEN_24184); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24785 = 6'hd == state ? $signed(w_4) : $signed(_GEN_24185); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24786 = 6'hd == state ? $signed(w_5) : $signed(_GEN_24186); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24787 = 6'hd == state ? $signed(w_6) : $signed(_GEN_24187); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24788 = 6'hd == state ? $signed(w_7) : $signed(_GEN_24188); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24789 = 6'hd == state ? $signed(w_8) : $signed(_GEN_24189); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24790 = 6'hd == state ? $signed(w_9) : $signed(_GEN_24190); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24791 = 6'hd == state ? $signed(w_10) : $signed(_GEN_24191); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24792 = 6'hd == state ? $signed(w_11) : $signed(_GEN_24192); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24793 = 6'hd == state ? $signed(w_12) : $signed(_GEN_24193); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24794 = 6'hd == state ? $signed(w_13) : $signed(_GEN_24194); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24795 = 6'hd == state ? $signed(w_14) : $signed(_GEN_24195); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24796 = 6'hd == state ? $signed(w_15) : $signed(_GEN_24196); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24797 = 6'hd == state ? $signed(w_16) : $signed(_GEN_24197); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24798 = 6'hd == state ? $signed(w_17) : $signed(_GEN_24198); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24799 = 6'hd == state ? $signed(w_18) : $signed(_GEN_24199); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24800 = 6'hd == state ? $signed(w_19) : $signed(_GEN_24200); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24801 = 6'hd == state ? $signed(w_20) : $signed(_GEN_24201); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24802 = 6'hd == state ? $signed(w_21) : $signed(_GEN_24202); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24803 = 6'hd == state ? $signed(w_22) : $signed(_GEN_24203); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24804 = 6'hd == state ? $signed(w_23) : $signed(_GEN_24204); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24805 = 6'hd == state ? $signed(w_24) : $signed(_GEN_24205); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24806 = 6'hd == state ? $signed(w_25) : $signed(_GEN_24206); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24807 = 6'hd == state ? $signed(w_26) : $signed(_GEN_24207); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24808 = 6'hd == state ? $signed(w_27) : $signed(_GEN_24208); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24809 = 6'hd == state ? $signed(w_28) : $signed(_GEN_24209); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24810 = 6'hd == state ? $signed(w_29) : $signed(_GEN_24210); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24811 = 6'hd == state ? $signed(w_30) : $signed(_GEN_24211); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24812 = 6'hd == state ? $signed(w_31) : $signed(_GEN_24212); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24813 = 6'hd == state ? $signed(w_32) : $signed(_GEN_24213); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24814 = 6'hd == state ? $signed(w_33) : $signed(_GEN_24214); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24815 = 6'hd == state ? $signed(w_34) : $signed(_GEN_24215); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24816 = 6'hd == state ? $signed(w_35) : $signed(_GEN_24216); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24817 = 6'hd == state ? $signed(w_36) : $signed(_GEN_24217); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24818 = 6'hd == state ? $signed(w_37) : $signed(_GEN_24218); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24819 = 6'hd == state ? $signed(w_38) : $signed(_GEN_24219); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24820 = 6'hd == state ? $signed(w_39) : $signed(_GEN_24220); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24821 = 6'hd == state ? $signed(w_40) : $signed(_GEN_24221); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24822 = 6'hd == state ? $signed(w_41) : $signed(_GEN_24222); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24823 = 6'hd == state ? $signed(w_42) : $signed(_GEN_24223); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24824 = 6'hd == state ? $signed(w_43) : $signed(_GEN_24224); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24825 = 6'hd == state ? $signed(w_44) : $signed(_GEN_24225); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24826 = 6'hd == state ? $signed(w_45) : $signed(_GEN_24226); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24827 = 6'hd == state ? $signed(w_46) : $signed(_GEN_24227); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24828 = 6'hd == state ? $signed(w_47) : $signed(_GEN_24228); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24829 = 6'hd == state ? $signed(w_48) : $signed(_GEN_24229); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24830 = 6'hd == state ? $signed(w_49) : $signed(_GEN_24230); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24831 = 6'hd == state ? $signed(w_50) : $signed(_GEN_24231); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24832 = 6'hd == state ? $signed(w_51) : $signed(_GEN_24232); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24833 = 6'hd == state ? $signed(w_52) : $signed(_GEN_24233); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24834 = 6'hd == state ? $signed(w_53) : $signed(_GEN_24234); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24835 = 6'hd == state ? $signed(w_54) : $signed(_GEN_24235); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24836 = 6'hd == state ? $signed(w_55) : $signed(_GEN_24236); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24837 = 6'hd == state ? $signed(w_56) : $signed(_GEN_24237); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24838 = 6'hd == state ? $signed(w_57) : $signed(_GEN_24238); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24839 = 6'hd == state ? $signed(w_58) : $signed(_GEN_24239); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24840 = 6'hd == state ? $signed(w_59) : $signed(_GEN_24240); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24841 = 6'hd == state ? $signed(w_60) : $signed(_GEN_24241); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24842 = 6'hd == state ? $signed(w_61) : $signed(_GEN_24242); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24843 = 6'hd == state ? $signed(w_62) : $signed(_GEN_24243); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24844 = 6'hd == state ? $signed(w_63) : $signed(_GEN_24244); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24845 = 6'hd == state ? $signed(w_64) : $signed(_GEN_24245); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24846 = 6'hd == state ? $signed(w_65) : $signed(_GEN_24246); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24847 = 6'hd == state ? $signed(w_66) : $signed(_GEN_24247); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24848 = 6'hd == state ? $signed(w_67) : $signed(_GEN_24248); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24849 = 6'hd == state ? $signed(w_68) : $signed(_GEN_24249); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24850 = 6'hd == state ? $signed(w_69) : $signed(_GEN_24250); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24851 = 6'hd == state ? $signed(w_70) : $signed(_GEN_24251); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24852 = 6'hd == state ? $signed(w_71) : $signed(_GEN_24252); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24853 = 6'hd == state ? $signed(w_72) : $signed(_GEN_24253); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24854 = 6'hd == state ? $signed(w_73) : $signed(_GEN_24254); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24855 = 6'hd == state ? $signed(w_74) : $signed(_GEN_24255); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24856 = 6'hd == state ? $signed(w_75) : $signed(_GEN_24256); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24857 = 6'hd == state ? $signed(w_76) : $signed(_GEN_24257); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24858 = 6'hd == state ? $signed(w_77) : $signed(_GEN_24258); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24859 = 6'hd == state ? $signed(w_78) : $signed(_GEN_24259); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24860 = 6'hd == state ? $signed(w_79) : $signed(_GEN_24260); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_24861 = 6'hd == state ? $signed(temp) : $signed(_GEN_24261); // @[digest.scala 38:19 81:19]
  wire  _GEN_24862 = 6'hd == state ? 1'h0 : _GEN_24262; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_24865 = 6'hd == state ? $signed(t) : $signed(_GEN_24265); // @[digest.scala 35:16 81:19]
  wire  _GEN_24866 = 6'hd == state ? 1'h0 : _GEN_24266; // @[digest.scala 81:19 48:24]
  wire [31:0] _GEN_24869 = 6'hd == state ? $signed(c) : $signed(_GEN_24270); // @[digest.scala 26:16 81:19]
  wire  _GEN_24870 = 6'hd == state ? 1'h0 : _GEN_24271; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_24873 = 6'hd == state ? $signed(b) : $signed(_GEN_24274); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_24874 = 6'hd == state ? $signed(a) : $signed(_GEN_24275); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_24956 = 6'hd == state ? $signed(digest_0) : $signed(_GEN_24357); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24957 = 6'hd == state ? $signed(digest_1) : $signed(_GEN_24358); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24958 = 6'hd == state ? $signed(digest_2) : $signed(_GEN_24359); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24959 = 6'hd == state ? $signed(digest_3) : $signed(_GEN_24360); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24960 = 6'hd == state ? $signed(digest_4) : $signed(_GEN_24361); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24961 = 6'hd == state ? $signed(digest_5) : $signed(_GEN_24362); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24962 = 6'hd == state ? $signed(digest_6) : $signed(_GEN_24363); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24963 = 6'hd == state ? $signed(digest_7) : $signed(_GEN_24364); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24964 = 6'hd == state ? $signed(digest_8) : $signed(_GEN_24365); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24965 = 6'hd == state ? $signed(digest_9) : $signed(_GEN_24366); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24966 = 6'hd == state ? $signed(digest_10) : $signed(_GEN_24367); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24967 = 6'hd == state ? $signed(digest_11) : $signed(_GEN_24368); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24968 = 6'hd == state ? $signed(digest_12) : $signed(_GEN_24369); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24969 = 6'hd == state ? $signed(digest_13) : $signed(_GEN_24370); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24970 = 6'hd == state ? $signed(digest_14) : $signed(_GEN_24371); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24971 = 6'hd == state ? $signed(digest_15) : $signed(_GEN_24372); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24972 = 6'hd == state ? $signed(digest_16) : $signed(_GEN_24373); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24973 = 6'hd == state ? $signed(digest_17) : $signed(_GEN_24374); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24974 = 6'hd == state ? $signed(digest_18) : $signed(_GEN_24375); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24975 = 6'hd == state ? $signed(digest_19) : $signed(_GEN_24376); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24976 = 6'hd == state ? $signed(digest_20) : $signed(_GEN_24377); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24977 = 6'hd == state ? $signed(digest_21) : $signed(_GEN_24378); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24978 = 6'hd == state ? $signed(digest_22) : $signed(_GEN_24379); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24979 = 6'hd == state ? $signed(digest_23) : $signed(_GEN_24380); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24980 = 6'hd == state ? $signed(digest_24) : $signed(_GEN_24381); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24981 = 6'hd == state ? $signed(digest_25) : $signed(_GEN_24382); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24982 = 6'hd == state ? $signed(digest_26) : $signed(_GEN_24383); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24983 = 6'hd == state ? $signed(digest_27) : $signed(_GEN_24384); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24984 = 6'hd == state ? $signed(digest_28) : $signed(_GEN_24385); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24985 = 6'hd == state ? $signed(digest_29) : $signed(_GEN_24386); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24986 = 6'hd == state ? $signed(digest_30) : $signed(_GEN_24387); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24987 = 6'hd == state ? $signed(digest_31) : $signed(_GEN_24388); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24988 = 6'hd == state ? $signed(digest_32) : $signed(_GEN_24389); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24989 = 6'hd == state ? $signed(digest_33) : $signed(_GEN_24390); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24990 = 6'hd == state ? $signed(digest_34) : $signed(_GEN_24391); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24991 = 6'hd == state ? $signed(digest_35) : $signed(_GEN_24392); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24992 = 6'hd == state ? $signed(digest_36) : $signed(_GEN_24393); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24993 = 6'hd == state ? $signed(digest_37) : $signed(_GEN_24394); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24994 = 6'hd == state ? $signed(digest_38) : $signed(_GEN_24395); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24995 = 6'hd == state ? $signed(digest_39) : $signed(_GEN_24396); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24996 = 6'hd == state ? $signed(digest_40) : $signed(_GEN_24397); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24997 = 6'hd == state ? $signed(digest_41) : $signed(_GEN_24398); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24998 = 6'hd == state ? $signed(digest_42) : $signed(_GEN_24399); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_24999 = 6'hd == state ? $signed(digest_43) : $signed(_GEN_24400); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25000 = 6'hd == state ? $signed(digest_44) : $signed(_GEN_24401); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25001 = 6'hd == state ? $signed(digest_45) : $signed(_GEN_24402); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25002 = 6'hd == state ? $signed(digest_46) : $signed(_GEN_24403); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25003 = 6'hd == state ? $signed(digest_47) : $signed(_GEN_24404); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25004 = 6'hd == state ? $signed(digest_48) : $signed(_GEN_24405); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25005 = 6'hd == state ? $signed(digest_49) : $signed(_GEN_24406); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25006 = 6'hd == state ? $signed(digest_50) : $signed(_GEN_24407); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25007 = 6'hd == state ? $signed(digest_51) : $signed(_GEN_24408); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25008 = 6'hd == state ? $signed(digest_52) : $signed(_GEN_24409); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25009 = 6'hd == state ? $signed(digest_53) : $signed(_GEN_24410); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25010 = 6'hd == state ? $signed(digest_54) : $signed(_GEN_24411); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25011 = 6'hd == state ? $signed(digest_55) : $signed(_GEN_24412); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25012 = 6'hd == state ? $signed(digest_56) : $signed(_GEN_24413); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25013 = 6'hd == state ? $signed(digest_57) : $signed(_GEN_24414); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25014 = 6'hd == state ? $signed(digest_58) : $signed(_GEN_24415); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25015 = 6'hd == state ? $signed(digest_59) : $signed(_GEN_24416); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25016 = 6'hd == state ? $signed(digest_60) : $signed(_GEN_24417); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25017 = 6'hd == state ? $signed(digest_61) : $signed(_GEN_24418); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25018 = 6'hd == state ? $signed(digest_62) : $signed(_GEN_24419); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25019 = 6'hd == state ? $signed(digest_63) : $signed(_GEN_24420); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25020 = 6'hd == state ? $signed(digest_64) : $signed(_GEN_24421); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25021 = 6'hd == state ? $signed(digest_65) : $signed(_GEN_24422); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25022 = 6'hd == state ? $signed(digest_66) : $signed(_GEN_24423); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25023 = 6'hd == state ? $signed(digest_67) : $signed(_GEN_24424); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25024 = 6'hd == state ? $signed(digest_68) : $signed(_GEN_24425); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25025 = 6'hd == state ? $signed(digest_69) : $signed(_GEN_24426); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25026 = 6'hd == state ? $signed(digest_70) : $signed(_GEN_24427); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25027 = 6'hd == state ? $signed(digest_71) : $signed(_GEN_24428); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25028 = 6'hd == state ? $signed(digest_72) : $signed(_GEN_24429); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25029 = 6'hd == state ? $signed(digest_73) : $signed(_GEN_24430); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25030 = 6'hd == state ? $signed(digest_74) : $signed(_GEN_24431); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25031 = 6'hd == state ? $signed(digest_75) : $signed(_GEN_24432); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25032 = 6'hd == state ? $signed(digest_76) : $signed(_GEN_24433); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25033 = 6'hd == state ? $signed(digest_77) : $signed(_GEN_24434); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25034 = 6'hd == state ? $signed(digest_78) : $signed(_GEN_24435); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25035 = 6'hd == state ? $signed(digest_79) : $signed(_GEN_24436); // @[digest.scala 81:19 53:21]
  wire  _GEN_25037 = 6'hd == state ? 1'h0 : _GEN_24438; // @[digest.scala 81:19 58:25]
  wire  _GEN_25120 = 6'hd == state ? 1'h0 : _GEN_24521; // @[digest.scala 81:19 63:25]
  wire  _GEN_25203 = 6'hd == state ? 1'h0 : _GEN_24604; // @[digest.scala 81:19 68:25]
  wire  _GEN_25286 = 6'hd == state ? 1'h0 : _GEN_24687; // @[digest.scala 81:19 73:25]
  wire  _GEN_25369 = 6'hd == state ? 1'h0 : _GEN_24770; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_25370 = 6'hc == state ? $signed(-32'sh67452302) : $signed(_GEN_24869); // @[digest.scala 133:15 81:19]
  wire [5:0] _GEN_25371 = 6'hc == state ? 6'hd : _GEN_24772; // @[digest.scala 134:19 81:19]
  wire [31:0] _GEN_25372 = 6'hc == state ? $signed(d) : $signed(_GEN_24771); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_25373 = 6'hc == state ? $signed(e) : $signed(_GEN_24773); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_25374 = 6'hc == state ? $signed(i) : $signed(_GEN_24774); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_25375 = 6'hc == state ? $signed(olda) : $signed(_GEN_24775); // @[digest.scala 29:19 81:19]
  wire [31:0] _GEN_25376 = 6'hc == state ? $signed(oldb) : $signed(_GEN_24776); // @[digest.scala 30:19 81:19]
  wire [31:0] _GEN_25377 = 6'hc == state ? $signed(oldc) : $signed(_GEN_24777); // @[digest.scala 31:19 81:19]
  wire [31:0] _GEN_25378 = 6'hc == state ? $signed(oldd) : $signed(_GEN_24778); // @[digest.scala 32:19 81:19]
  wire [31:0] _GEN_25379 = 6'hc == state ? $signed(olde) : $signed(_GEN_24779); // @[digest.scala 33:19 81:19]
  wire [31:0] _GEN_25380 = 6'hc == state ? $signed(j) : $signed(_GEN_24780); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_25381 = 6'hc == state ? $signed(w_0) : $signed(_GEN_24781); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25382 = 6'hc == state ? $signed(w_1) : $signed(_GEN_24782); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25383 = 6'hc == state ? $signed(w_2) : $signed(_GEN_24783); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25384 = 6'hc == state ? $signed(w_3) : $signed(_GEN_24784); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25385 = 6'hc == state ? $signed(w_4) : $signed(_GEN_24785); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25386 = 6'hc == state ? $signed(w_5) : $signed(_GEN_24786); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25387 = 6'hc == state ? $signed(w_6) : $signed(_GEN_24787); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25388 = 6'hc == state ? $signed(w_7) : $signed(_GEN_24788); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25389 = 6'hc == state ? $signed(w_8) : $signed(_GEN_24789); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25390 = 6'hc == state ? $signed(w_9) : $signed(_GEN_24790); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25391 = 6'hc == state ? $signed(w_10) : $signed(_GEN_24791); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25392 = 6'hc == state ? $signed(w_11) : $signed(_GEN_24792); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25393 = 6'hc == state ? $signed(w_12) : $signed(_GEN_24793); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25394 = 6'hc == state ? $signed(w_13) : $signed(_GEN_24794); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25395 = 6'hc == state ? $signed(w_14) : $signed(_GEN_24795); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25396 = 6'hc == state ? $signed(w_15) : $signed(_GEN_24796); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25397 = 6'hc == state ? $signed(w_16) : $signed(_GEN_24797); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25398 = 6'hc == state ? $signed(w_17) : $signed(_GEN_24798); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25399 = 6'hc == state ? $signed(w_18) : $signed(_GEN_24799); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25400 = 6'hc == state ? $signed(w_19) : $signed(_GEN_24800); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25401 = 6'hc == state ? $signed(w_20) : $signed(_GEN_24801); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25402 = 6'hc == state ? $signed(w_21) : $signed(_GEN_24802); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25403 = 6'hc == state ? $signed(w_22) : $signed(_GEN_24803); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25404 = 6'hc == state ? $signed(w_23) : $signed(_GEN_24804); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25405 = 6'hc == state ? $signed(w_24) : $signed(_GEN_24805); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25406 = 6'hc == state ? $signed(w_25) : $signed(_GEN_24806); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25407 = 6'hc == state ? $signed(w_26) : $signed(_GEN_24807); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25408 = 6'hc == state ? $signed(w_27) : $signed(_GEN_24808); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25409 = 6'hc == state ? $signed(w_28) : $signed(_GEN_24809); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25410 = 6'hc == state ? $signed(w_29) : $signed(_GEN_24810); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25411 = 6'hc == state ? $signed(w_30) : $signed(_GEN_24811); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25412 = 6'hc == state ? $signed(w_31) : $signed(_GEN_24812); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25413 = 6'hc == state ? $signed(w_32) : $signed(_GEN_24813); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25414 = 6'hc == state ? $signed(w_33) : $signed(_GEN_24814); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25415 = 6'hc == state ? $signed(w_34) : $signed(_GEN_24815); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25416 = 6'hc == state ? $signed(w_35) : $signed(_GEN_24816); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25417 = 6'hc == state ? $signed(w_36) : $signed(_GEN_24817); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25418 = 6'hc == state ? $signed(w_37) : $signed(_GEN_24818); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25419 = 6'hc == state ? $signed(w_38) : $signed(_GEN_24819); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25420 = 6'hc == state ? $signed(w_39) : $signed(_GEN_24820); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25421 = 6'hc == state ? $signed(w_40) : $signed(_GEN_24821); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25422 = 6'hc == state ? $signed(w_41) : $signed(_GEN_24822); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25423 = 6'hc == state ? $signed(w_42) : $signed(_GEN_24823); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25424 = 6'hc == state ? $signed(w_43) : $signed(_GEN_24824); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25425 = 6'hc == state ? $signed(w_44) : $signed(_GEN_24825); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25426 = 6'hc == state ? $signed(w_45) : $signed(_GEN_24826); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25427 = 6'hc == state ? $signed(w_46) : $signed(_GEN_24827); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25428 = 6'hc == state ? $signed(w_47) : $signed(_GEN_24828); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25429 = 6'hc == state ? $signed(w_48) : $signed(_GEN_24829); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25430 = 6'hc == state ? $signed(w_49) : $signed(_GEN_24830); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25431 = 6'hc == state ? $signed(w_50) : $signed(_GEN_24831); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25432 = 6'hc == state ? $signed(w_51) : $signed(_GEN_24832); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25433 = 6'hc == state ? $signed(w_52) : $signed(_GEN_24833); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25434 = 6'hc == state ? $signed(w_53) : $signed(_GEN_24834); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25435 = 6'hc == state ? $signed(w_54) : $signed(_GEN_24835); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25436 = 6'hc == state ? $signed(w_55) : $signed(_GEN_24836); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25437 = 6'hc == state ? $signed(w_56) : $signed(_GEN_24837); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25438 = 6'hc == state ? $signed(w_57) : $signed(_GEN_24838); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25439 = 6'hc == state ? $signed(w_58) : $signed(_GEN_24839); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25440 = 6'hc == state ? $signed(w_59) : $signed(_GEN_24840); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25441 = 6'hc == state ? $signed(w_60) : $signed(_GEN_24841); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25442 = 6'hc == state ? $signed(w_61) : $signed(_GEN_24842); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25443 = 6'hc == state ? $signed(w_62) : $signed(_GEN_24843); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25444 = 6'hc == state ? $signed(w_63) : $signed(_GEN_24844); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25445 = 6'hc == state ? $signed(w_64) : $signed(_GEN_24845); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25446 = 6'hc == state ? $signed(w_65) : $signed(_GEN_24846); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25447 = 6'hc == state ? $signed(w_66) : $signed(_GEN_24847); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25448 = 6'hc == state ? $signed(w_67) : $signed(_GEN_24848); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25449 = 6'hc == state ? $signed(w_68) : $signed(_GEN_24849); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25450 = 6'hc == state ? $signed(w_69) : $signed(_GEN_24850); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25451 = 6'hc == state ? $signed(w_70) : $signed(_GEN_24851); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25452 = 6'hc == state ? $signed(w_71) : $signed(_GEN_24852); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25453 = 6'hc == state ? $signed(w_72) : $signed(_GEN_24853); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25454 = 6'hc == state ? $signed(w_73) : $signed(_GEN_24854); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25455 = 6'hc == state ? $signed(w_74) : $signed(_GEN_24855); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25456 = 6'hc == state ? $signed(w_75) : $signed(_GEN_24856); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25457 = 6'hc == state ? $signed(w_76) : $signed(_GEN_24857); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25458 = 6'hc == state ? $signed(w_77) : $signed(_GEN_24858); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25459 = 6'hc == state ? $signed(w_78) : $signed(_GEN_24859); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25460 = 6'hc == state ? $signed(w_79) : $signed(_GEN_24860); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25461 = 6'hc == state ? $signed(temp) : $signed(_GEN_24861); // @[digest.scala 38:19 81:19]
  wire  _GEN_25462 = 6'hc == state ? 1'h0 : _GEN_24862; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_25465 = 6'hc == state ? $signed(t) : $signed(_GEN_24865); // @[digest.scala 35:16 81:19]
  wire  _GEN_25466 = 6'hc == state ? 1'h0 : _GEN_24866; // @[digest.scala 81:19 48:24]
  wire  _GEN_25469 = 6'hc == state ? 1'h0 : _GEN_24870; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_25472 = 6'hc == state ? $signed(b) : $signed(_GEN_24873); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_25473 = 6'hc == state ? $signed(a) : $signed(_GEN_24874); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_25555 = 6'hc == state ? $signed(digest_0) : $signed(_GEN_24956); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25556 = 6'hc == state ? $signed(digest_1) : $signed(_GEN_24957); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25557 = 6'hc == state ? $signed(digest_2) : $signed(_GEN_24958); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25558 = 6'hc == state ? $signed(digest_3) : $signed(_GEN_24959); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25559 = 6'hc == state ? $signed(digest_4) : $signed(_GEN_24960); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25560 = 6'hc == state ? $signed(digest_5) : $signed(_GEN_24961); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25561 = 6'hc == state ? $signed(digest_6) : $signed(_GEN_24962); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25562 = 6'hc == state ? $signed(digest_7) : $signed(_GEN_24963); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25563 = 6'hc == state ? $signed(digest_8) : $signed(_GEN_24964); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25564 = 6'hc == state ? $signed(digest_9) : $signed(_GEN_24965); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25565 = 6'hc == state ? $signed(digest_10) : $signed(_GEN_24966); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25566 = 6'hc == state ? $signed(digest_11) : $signed(_GEN_24967); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25567 = 6'hc == state ? $signed(digest_12) : $signed(_GEN_24968); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25568 = 6'hc == state ? $signed(digest_13) : $signed(_GEN_24969); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25569 = 6'hc == state ? $signed(digest_14) : $signed(_GEN_24970); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25570 = 6'hc == state ? $signed(digest_15) : $signed(_GEN_24971); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25571 = 6'hc == state ? $signed(digest_16) : $signed(_GEN_24972); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25572 = 6'hc == state ? $signed(digest_17) : $signed(_GEN_24973); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25573 = 6'hc == state ? $signed(digest_18) : $signed(_GEN_24974); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25574 = 6'hc == state ? $signed(digest_19) : $signed(_GEN_24975); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25575 = 6'hc == state ? $signed(digest_20) : $signed(_GEN_24976); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25576 = 6'hc == state ? $signed(digest_21) : $signed(_GEN_24977); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25577 = 6'hc == state ? $signed(digest_22) : $signed(_GEN_24978); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25578 = 6'hc == state ? $signed(digest_23) : $signed(_GEN_24979); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25579 = 6'hc == state ? $signed(digest_24) : $signed(_GEN_24980); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25580 = 6'hc == state ? $signed(digest_25) : $signed(_GEN_24981); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25581 = 6'hc == state ? $signed(digest_26) : $signed(_GEN_24982); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25582 = 6'hc == state ? $signed(digest_27) : $signed(_GEN_24983); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25583 = 6'hc == state ? $signed(digest_28) : $signed(_GEN_24984); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25584 = 6'hc == state ? $signed(digest_29) : $signed(_GEN_24985); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25585 = 6'hc == state ? $signed(digest_30) : $signed(_GEN_24986); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25586 = 6'hc == state ? $signed(digest_31) : $signed(_GEN_24987); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25587 = 6'hc == state ? $signed(digest_32) : $signed(_GEN_24988); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25588 = 6'hc == state ? $signed(digest_33) : $signed(_GEN_24989); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25589 = 6'hc == state ? $signed(digest_34) : $signed(_GEN_24990); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25590 = 6'hc == state ? $signed(digest_35) : $signed(_GEN_24991); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25591 = 6'hc == state ? $signed(digest_36) : $signed(_GEN_24992); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25592 = 6'hc == state ? $signed(digest_37) : $signed(_GEN_24993); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25593 = 6'hc == state ? $signed(digest_38) : $signed(_GEN_24994); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25594 = 6'hc == state ? $signed(digest_39) : $signed(_GEN_24995); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25595 = 6'hc == state ? $signed(digest_40) : $signed(_GEN_24996); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25596 = 6'hc == state ? $signed(digest_41) : $signed(_GEN_24997); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25597 = 6'hc == state ? $signed(digest_42) : $signed(_GEN_24998); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25598 = 6'hc == state ? $signed(digest_43) : $signed(_GEN_24999); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25599 = 6'hc == state ? $signed(digest_44) : $signed(_GEN_25000); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25600 = 6'hc == state ? $signed(digest_45) : $signed(_GEN_25001); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25601 = 6'hc == state ? $signed(digest_46) : $signed(_GEN_25002); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25602 = 6'hc == state ? $signed(digest_47) : $signed(_GEN_25003); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25603 = 6'hc == state ? $signed(digest_48) : $signed(_GEN_25004); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25604 = 6'hc == state ? $signed(digest_49) : $signed(_GEN_25005); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25605 = 6'hc == state ? $signed(digest_50) : $signed(_GEN_25006); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25606 = 6'hc == state ? $signed(digest_51) : $signed(_GEN_25007); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25607 = 6'hc == state ? $signed(digest_52) : $signed(_GEN_25008); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25608 = 6'hc == state ? $signed(digest_53) : $signed(_GEN_25009); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25609 = 6'hc == state ? $signed(digest_54) : $signed(_GEN_25010); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25610 = 6'hc == state ? $signed(digest_55) : $signed(_GEN_25011); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25611 = 6'hc == state ? $signed(digest_56) : $signed(_GEN_25012); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25612 = 6'hc == state ? $signed(digest_57) : $signed(_GEN_25013); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25613 = 6'hc == state ? $signed(digest_58) : $signed(_GEN_25014); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25614 = 6'hc == state ? $signed(digest_59) : $signed(_GEN_25015); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25615 = 6'hc == state ? $signed(digest_60) : $signed(_GEN_25016); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25616 = 6'hc == state ? $signed(digest_61) : $signed(_GEN_25017); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25617 = 6'hc == state ? $signed(digest_62) : $signed(_GEN_25018); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25618 = 6'hc == state ? $signed(digest_63) : $signed(_GEN_25019); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25619 = 6'hc == state ? $signed(digest_64) : $signed(_GEN_25020); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25620 = 6'hc == state ? $signed(digest_65) : $signed(_GEN_25021); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25621 = 6'hc == state ? $signed(digest_66) : $signed(_GEN_25022); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25622 = 6'hc == state ? $signed(digest_67) : $signed(_GEN_25023); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25623 = 6'hc == state ? $signed(digest_68) : $signed(_GEN_25024); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25624 = 6'hc == state ? $signed(digest_69) : $signed(_GEN_25025); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25625 = 6'hc == state ? $signed(digest_70) : $signed(_GEN_25026); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25626 = 6'hc == state ? $signed(digest_71) : $signed(_GEN_25027); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25627 = 6'hc == state ? $signed(digest_72) : $signed(_GEN_25028); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25628 = 6'hc == state ? $signed(digest_73) : $signed(_GEN_25029); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25629 = 6'hc == state ? $signed(digest_74) : $signed(_GEN_25030); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25630 = 6'hc == state ? $signed(digest_75) : $signed(_GEN_25031); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25631 = 6'hc == state ? $signed(digest_76) : $signed(_GEN_25032); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25632 = 6'hc == state ? $signed(digest_77) : $signed(_GEN_25033); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25633 = 6'hc == state ? $signed(digest_78) : $signed(_GEN_25034); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_25634 = 6'hc == state ? $signed(digest_79) : $signed(_GEN_25035); // @[digest.scala 81:19 53:21]
  wire  _GEN_25636 = 6'hc == state ? 1'h0 : _GEN_25037; // @[digest.scala 81:19 58:25]
  wire  _GEN_25719 = 6'hc == state ? 1'h0 : _GEN_25120; // @[digest.scala 81:19 63:25]
  wire  _GEN_25802 = 6'hc == state ? 1'h0 : _GEN_25203; // @[digest.scala 81:19 68:25]
  wire  _GEN_25885 = 6'hc == state ? 1'h0 : _GEN_25286; // @[digest.scala 81:19 73:25]
  wire  _GEN_25968 = 6'hc == state ? 1'h0 : _GEN_25369; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_25969 = 6'hb == state ? $signed(-32'sh10325477) : $signed(_GEN_25472); // @[digest.scala 129:15 81:19]
  wire [5:0] _GEN_25970 = 6'hb == state ? 6'hc : _GEN_25371; // @[digest.scala 130:19 81:19]
  wire [31:0] _GEN_25971 = 6'hb == state ? $signed(c) : $signed(_GEN_25370); // @[digest.scala 26:16 81:19]
  wire [31:0] _GEN_25972 = 6'hb == state ? $signed(d) : $signed(_GEN_25372); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_25973 = 6'hb == state ? $signed(e) : $signed(_GEN_25373); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_25974 = 6'hb == state ? $signed(i) : $signed(_GEN_25374); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_25975 = 6'hb == state ? $signed(olda) : $signed(_GEN_25375); // @[digest.scala 29:19 81:19]
  wire [31:0] _GEN_25976 = 6'hb == state ? $signed(oldb) : $signed(_GEN_25376); // @[digest.scala 30:19 81:19]
  wire [31:0] _GEN_25977 = 6'hb == state ? $signed(oldc) : $signed(_GEN_25377); // @[digest.scala 31:19 81:19]
  wire [31:0] _GEN_25978 = 6'hb == state ? $signed(oldd) : $signed(_GEN_25378); // @[digest.scala 32:19 81:19]
  wire [31:0] _GEN_25979 = 6'hb == state ? $signed(olde) : $signed(_GEN_25379); // @[digest.scala 33:19 81:19]
  wire [31:0] _GEN_25980 = 6'hb == state ? $signed(j) : $signed(_GEN_25380); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_25981 = 6'hb == state ? $signed(w_0) : $signed(_GEN_25381); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25982 = 6'hb == state ? $signed(w_1) : $signed(_GEN_25382); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25983 = 6'hb == state ? $signed(w_2) : $signed(_GEN_25383); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25984 = 6'hb == state ? $signed(w_3) : $signed(_GEN_25384); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25985 = 6'hb == state ? $signed(w_4) : $signed(_GEN_25385); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25986 = 6'hb == state ? $signed(w_5) : $signed(_GEN_25386); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25987 = 6'hb == state ? $signed(w_6) : $signed(_GEN_25387); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25988 = 6'hb == state ? $signed(w_7) : $signed(_GEN_25388); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25989 = 6'hb == state ? $signed(w_8) : $signed(_GEN_25389); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25990 = 6'hb == state ? $signed(w_9) : $signed(_GEN_25390); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25991 = 6'hb == state ? $signed(w_10) : $signed(_GEN_25391); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25992 = 6'hb == state ? $signed(w_11) : $signed(_GEN_25392); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25993 = 6'hb == state ? $signed(w_12) : $signed(_GEN_25393); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25994 = 6'hb == state ? $signed(w_13) : $signed(_GEN_25394); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25995 = 6'hb == state ? $signed(w_14) : $signed(_GEN_25395); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25996 = 6'hb == state ? $signed(w_15) : $signed(_GEN_25396); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25997 = 6'hb == state ? $signed(w_16) : $signed(_GEN_25397); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25998 = 6'hb == state ? $signed(w_17) : $signed(_GEN_25398); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_25999 = 6'hb == state ? $signed(w_18) : $signed(_GEN_25399); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26000 = 6'hb == state ? $signed(w_19) : $signed(_GEN_25400); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26001 = 6'hb == state ? $signed(w_20) : $signed(_GEN_25401); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26002 = 6'hb == state ? $signed(w_21) : $signed(_GEN_25402); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26003 = 6'hb == state ? $signed(w_22) : $signed(_GEN_25403); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26004 = 6'hb == state ? $signed(w_23) : $signed(_GEN_25404); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26005 = 6'hb == state ? $signed(w_24) : $signed(_GEN_25405); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26006 = 6'hb == state ? $signed(w_25) : $signed(_GEN_25406); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26007 = 6'hb == state ? $signed(w_26) : $signed(_GEN_25407); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26008 = 6'hb == state ? $signed(w_27) : $signed(_GEN_25408); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26009 = 6'hb == state ? $signed(w_28) : $signed(_GEN_25409); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26010 = 6'hb == state ? $signed(w_29) : $signed(_GEN_25410); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26011 = 6'hb == state ? $signed(w_30) : $signed(_GEN_25411); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26012 = 6'hb == state ? $signed(w_31) : $signed(_GEN_25412); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26013 = 6'hb == state ? $signed(w_32) : $signed(_GEN_25413); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26014 = 6'hb == state ? $signed(w_33) : $signed(_GEN_25414); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26015 = 6'hb == state ? $signed(w_34) : $signed(_GEN_25415); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26016 = 6'hb == state ? $signed(w_35) : $signed(_GEN_25416); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26017 = 6'hb == state ? $signed(w_36) : $signed(_GEN_25417); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26018 = 6'hb == state ? $signed(w_37) : $signed(_GEN_25418); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26019 = 6'hb == state ? $signed(w_38) : $signed(_GEN_25419); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26020 = 6'hb == state ? $signed(w_39) : $signed(_GEN_25420); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26021 = 6'hb == state ? $signed(w_40) : $signed(_GEN_25421); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26022 = 6'hb == state ? $signed(w_41) : $signed(_GEN_25422); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26023 = 6'hb == state ? $signed(w_42) : $signed(_GEN_25423); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26024 = 6'hb == state ? $signed(w_43) : $signed(_GEN_25424); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26025 = 6'hb == state ? $signed(w_44) : $signed(_GEN_25425); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26026 = 6'hb == state ? $signed(w_45) : $signed(_GEN_25426); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26027 = 6'hb == state ? $signed(w_46) : $signed(_GEN_25427); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26028 = 6'hb == state ? $signed(w_47) : $signed(_GEN_25428); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26029 = 6'hb == state ? $signed(w_48) : $signed(_GEN_25429); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26030 = 6'hb == state ? $signed(w_49) : $signed(_GEN_25430); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26031 = 6'hb == state ? $signed(w_50) : $signed(_GEN_25431); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26032 = 6'hb == state ? $signed(w_51) : $signed(_GEN_25432); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26033 = 6'hb == state ? $signed(w_52) : $signed(_GEN_25433); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26034 = 6'hb == state ? $signed(w_53) : $signed(_GEN_25434); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26035 = 6'hb == state ? $signed(w_54) : $signed(_GEN_25435); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26036 = 6'hb == state ? $signed(w_55) : $signed(_GEN_25436); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26037 = 6'hb == state ? $signed(w_56) : $signed(_GEN_25437); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26038 = 6'hb == state ? $signed(w_57) : $signed(_GEN_25438); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26039 = 6'hb == state ? $signed(w_58) : $signed(_GEN_25439); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26040 = 6'hb == state ? $signed(w_59) : $signed(_GEN_25440); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26041 = 6'hb == state ? $signed(w_60) : $signed(_GEN_25441); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26042 = 6'hb == state ? $signed(w_61) : $signed(_GEN_25442); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26043 = 6'hb == state ? $signed(w_62) : $signed(_GEN_25443); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26044 = 6'hb == state ? $signed(w_63) : $signed(_GEN_25444); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26045 = 6'hb == state ? $signed(w_64) : $signed(_GEN_25445); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26046 = 6'hb == state ? $signed(w_65) : $signed(_GEN_25446); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26047 = 6'hb == state ? $signed(w_66) : $signed(_GEN_25447); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26048 = 6'hb == state ? $signed(w_67) : $signed(_GEN_25448); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26049 = 6'hb == state ? $signed(w_68) : $signed(_GEN_25449); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26050 = 6'hb == state ? $signed(w_69) : $signed(_GEN_25450); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26051 = 6'hb == state ? $signed(w_70) : $signed(_GEN_25451); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26052 = 6'hb == state ? $signed(w_71) : $signed(_GEN_25452); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26053 = 6'hb == state ? $signed(w_72) : $signed(_GEN_25453); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26054 = 6'hb == state ? $signed(w_73) : $signed(_GEN_25454); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26055 = 6'hb == state ? $signed(w_74) : $signed(_GEN_25455); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26056 = 6'hb == state ? $signed(w_75) : $signed(_GEN_25456); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26057 = 6'hb == state ? $signed(w_76) : $signed(_GEN_25457); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26058 = 6'hb == state ? $signed(w_77) : $signed(_GEN_25458); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26059 = 6'hb == state ? $signed(w_78) : $signed(_GEN_25459); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26060 = 6'hb == state ? $signed(w_79) : $signed(_GEN_25460); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26061 = 6'hb == state ? $signed(temp) : $signed(_GEN_25461); // @[digest.scala 38:19 81:19]
  wire  _GEN_26062 = 6'hb == state ? 1'h0 : _GEN_25462; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_26065 = 6'hb == state ? $signed(t) : $signed(_GEN_25465); // @[digest.scala 35:16 81:19]
  wire  _GEN_26066 = 6'hb == state ? 1'h0 : _GEN_25466; // @[digest.scala 81:19 48:24]
  wire  _GEN_26069 = 6'hb == state ? 1'h0 : _GEN_25469; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_26072 = 6'hb == state ? $signed(a) : $signed(_GEN_25473); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_26154 = 6'hb == state ? $signed(digest_0) : $signed(_GEN_25555); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26155 = 6'hb == state ? $signed(digest_1) : $signed(_GEN_25556); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26156 = 6'hb == state ? $signed(digest_2) : $signed(_GEN_25557); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26157 = 6'hb == state ? $signed(digest_3) : $signed(_GEN_25558); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26158 = 6'hb == state ? $signed(digest_4) : $signed(_GEN_25559); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26159 = 6'hb == state ? $signed(digest_5) : $signed(_GEN_25560); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26160 = 6'hb == state ? $signed(digest_6) : $signed(_GEN_25561); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26161 = 6'hb == state ? $signed(digest_7) : $signed(_GEN_25562); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26162 = 6'hb == state ? $signed(digest_8) : $signed(_GEN_25563); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26163 = 6'hb == state ? $signed(digest_9) : $signed(_GEN_25564); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26164 = 6'hb == state ? $signed(digest_10) : $signed(_GEN_25565); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26165 = 6'hb == state ? $signed(digest_11) : $signed(_GEN_25566); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26166 = 6'hb == state ? $signed(digest_12) : $signed(_GEN_25567); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26167 = 6'hb == state ? $signed(digest_13) : $signed(_GEN_25568); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26168 = 6'hb == state ? $signed(digest_14) : $signed(_GEN_25569); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26169 = 6'hb == state ? $signed(digest_15) : $signed(_GEN_25570); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26170 = 6'hb == state ? $signed(digest_16) : $signed(_GEN_25571); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26171 = 6'hb == state ? $signed(digest_17) : $signed(_GEN_25572); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26172 = 6'hb == state ? $signed(digest_18) : $signed(_GEN_25573); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26173 = 6'hb == state ? $signed(digest_19) : $signed(_GEN_25574); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26174 = 6'hb == state ? $signed(digest_20) : $signed(_GEN_25575); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26175 = 6'hb == state ? $signed(digest_21) : $signed(_GEN_25576); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26176 = 6'hb == state ? $signed(digest_22) : $signed(_GEN_25577); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26177 = 6'hb == state ? $signed(digest_23) : $signed(_GEN_25578); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26178 = 6'hb == state ? $signed(digest_24) : $signed(_GEN_25579); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26179 = 6'hb == state ? $signed(digest_25) : $signed(_GEN_25580); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26180 = 6'hb == state ? $signed(digest_26) : $signed(_GEN_25581); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26181 = 6'hb == state ? $signed(digest_27) : $signed(_GEN_25582); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26182 = 6'hb == state ? $signed(digest_28) : $signed(_GEN_25583); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26183 = 6'hb == state ? $signed(digest_29) : $signed(_GEN_25584); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26184 = 6'hb == state ? $signed(digest_30) : $signed(_GEN_25585); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26185 = 6'hb == state ? $signed(digest_31) : $signed(_GEN_25586); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26186 = 6'hb == state ? $signed(digest_32) : $signed(_GEN_25587); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26187 = 6'hb == state ? $signed(digest_33) : $signed(_GEN_25588); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26188 = 6'hb == state ? $signed(digest_34) : $signed(_GEN_25589); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26189 = 6'hb == state ? $signed(digest_35) : $signed(_GEN_25590); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26190 = 6'hb == state ? $signed(digest_36) : $signed(_GEN_25591); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26191 = 6'hb == state ? $signed(digest_37) : $signed(_GEN_25592); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26192 = 6'hb == state ? $signed(digest_38) : $signed(_GEN_25593); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26193 = 6'hb == state ? $signed(digest_39) : $signed(_GEN_25594); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26194 = 6'hb == state ? $signed(digest_40) : $signed(_GEN_25595); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26195 = 6'hb == state ? $signed(digest_41) : $signed(_GEN_25596); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26196 = 6'hb == state ? $signed(digest_42) : $signed(_GEN_25597); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26197 = 6'hb == state ? $signed(digest_43) : $signed(_GEN_25598); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26198 = 6'hb == state ? $signed(digest_44) : $signed(_GEN_25599); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26199 = 6'hb == state ? $signed(digest_45) : $signed(_GEN_25600); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26200 = 6'hb == state ? $signed(digest_46) : $signed(_GEN_25601); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26201 = 6'hb == state ? $signed(digest_47) : $signed(_GEN_25602); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26202 = 6'hb == state ? $signed(digest_48) : $signed(_GEN_25603); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26203 = 6'hb == state ? $signed(digest_49) : $signed(_GEN_25604); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26204 = 6'hb == state ? $signed(digest_50) : $signed(_GEN_25605); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26205 = 6'hb == state ? $signed(digest_51) : $signed(_GEN_25606); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26206 = 6'hb == state ? $signed(digest_52) : $signed(_GEN_25607); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26207 = 6'hb == state ? $signed(digest_53) : $signed(_GEN_25608); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26208 = 6'hb == state ? $signed(digest_54) : $signed(_GEN_25609); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26209 = 6'hb == state ? $signed(digest_55) : $signed(_GEN_25610); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26210 = 6'hb == state ? $signed(digest_56) : $signed(_GEN_25611); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26211 = 6'hb == state ? $signed(digest_57) : $signed(_GEN_25612); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26212 = 6'hb == state ? $signed(digest_58) : $signed(_GEN_25613); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26213 = 6'hb == state ? $signed(digest_59) : $signed(_GEN_25614); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26214 = 6'hb == state ? $signed(digest_60) : $signed(_GEN_25615); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26215 = 6'hb == state ? $signed(digest_61) : $signed(_GEN_25616); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26216 = 6'hb == state ? $signed(digest_62) : $signed(_GEN_25617); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26217 = 6'hb == state ? $signed(digest_63) : $signed(_GEN_25618); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26218 = 6'hb == state ? $signed(digest_64) : $signed(_GEN_25619); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26219 = 6'hb == state ? $signed(digest_65) : $signed(_GEN_25620); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26220 = 6'hb == state ? $signed(digest_66) : $signed(_GEN_25621); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26221 = 6'hb == state ? $signed(digest_67) : $signed(_GEN_25622); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26222 = 6'hb == state ? $signed(digest_68) : $signed(_GEN_25623); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26223 = 6'hb == state ? $signed(digest_69) : $signed(_GEN_25624); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26224 = 6'hb == state ? $signed(digest_70) : $signed(_GEN_25625); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26225 = 6'hb == state ? $signed(digest_71) : $signed(_GEN_25626); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26226 = 6'hb == state ? $signed(digest_72) : $signed(_GEN_25627); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26227 = 6'hb == state ? $signed(digest_73) : $signed(_GEN_25628); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26228 = 6'hb == state ? $signed(digest_74) : $signed(_GEN_25629); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26229 = 6'hb == state ? $signed(digest_75) : $signed(_GEN_25630); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26230 = 6'hb == state ? $signed(digest_76) : $signed(_GEN_25631); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26231 = 6'hb == state ? $signed(digest_77) : $signed(_GEN_25632); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26232 = 6'hb == state ? $signed(digest_78) : $signed(_GEN_25633); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26233 = 6'hb == state ? $signed(digest_79) : $signed(_GEN_25634); // @[digest.scala 81:19 53:21]
  wire  _GEN_26235 = 6'hb == state ? 1'h0 : _GEN_25636; // @[digest.scala 81:19 58:25]
  wire  _GEN_26318 = 6'hb == state ? 1'h0 : _GEN_25719; // @[digest.scala 81:19 63:25]
  wire  _GEN_26401 = 6'hb == state ? 1'h0 : _GEN_25802; // @[digest.scala 81:19 68:25]
  wire  _GEN_26484 = 6'hb == state ? 1'h0 : _GEN_25885; // @[digest.scala 81:19 73:25]
  wire  _GEN_26567 = 6'hb == state ? 1'h0 : _GEN_25968; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_26568 = 6'ha == state ? $signed(32'sh67452301) : $signed(_GEN_26072); // @[digest.scala 125:15 81:19]
  wire [5:0] _GEN_26569 = 6'ha == state ? 6'hb : _GEN_25970; // @[digest.scala 126:19 81:19]
  wire [31:0] _GEN_26570 = 6'ha == state ? $signed(b) : $signed(_GEN_25969); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_26571 = 6'ha == state ? $signed(c) : $signed(_GEN_25971); // @[digest.scala 26:16 81:19]
  wire [31:0] _GEN_26572 = 6'ha == state ? $signed(d) : $signed(_GEN_25972); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_26573 = 6'ha == state ? $signed(e) : $signed(_GEN_25973); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_26574 = 6'ha == state ? $signed(i) : $signed(_GEN_25974); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_26575 = 6'ha == state ? $signed(olda) : $signed(_GEN_25975); // @[digest.scala 29:19 81:19]
  wire [31:0] _GEN_26576 = 6'ha == state ? $signed(oldb) : $signed(_GEN_25976); // @[digest.scala 30:19 81:19]
  wire [31:0] _GEN_26577 = 6'ha == state ? $signed(oldc) : $signed(_GEN_25977); // @[digest.scala 31:19 81:19]
  wire [31:0] _GEN_26578 = 6'ha == state ? $signed(oldd) : $signed(_GEN_25978); // @[digest.scala 32:19 81:19]
  wire [31:0] _GEN_26579 = 6'ha == state ? $signed(olde) : $signed(_GEN_25979); // @[digest.scala 33:19 81:19]
  wire [31:0] _GEN_26580 = 6'ha == state ? $signed(j) : $signed(_GEN_25980); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_26581 = 6'ha == state ? $signed(w_0) : $signed(_GEN_25981); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26582 = 6'ha == state ? $signed(w_1) : $signed(_GEN_25982); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26583 = 6'ha == state ? $signed(w_2) : $signed(_GEN_25983); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26584 = 6'ha == state ? $signed(w_3) : $signed(_GEN_25984); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26585 = 6'ha == state ? $signed(w_4) : $signed(_GEN_25985); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26586 = 6'ha == state ? $signed(w_5) : $signed(_GEN_25986); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26587 = 6'ha == state ? $signed(w_6) : $signed(_GEN_25987); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26588 = 6'ha == state ? $signed(w_7) : $signed(_GEN_25988); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26589 = 6'ha == state ? $signed(w_8) : $signed(_GEN_25989); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26590 = 6'ha == state ? $signed(w_9) : $signed(_GEN_25990); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26591 = 6'ha == state ? $signed(w_10) : $signed(_GEN_25991); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26592 = 6'ha == state ? $signed(w_11) : $signed(_GEN_25992); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26593 = 6'ha == state ? $signed(w_12) : $signed(_GEN_25993); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26594 = 6'ha == state ? $signed(w_13) : $signed(_GEN_25994); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26595 = 6'ha == state ? $signed(w_14) : $signed(_GEN_25995); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26596 = 6'ha == state ? $signed(w_15) : $signed(_GEN_25996); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26597 = 6'ha == state ? $signed(w_16) : $signed(_GEN_25997); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26598 = 6'ha == state ? $signed(w_17) : $signed(_GEN_25998); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26599 = 6'ha == state ? $signed(w_18) : $signed(_GEN_25999); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26600 = 6'ha == state ? $signed(w_19) : $signed(_GEN_26000); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26601 = 6'ha == state ? $signed(w_20) : $signed(_GEN_26001); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26602 = 6'ha == state ? $signed(w_21) : $signed(_GEN_26002); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26603 = 6'ha == state ? $signed(w_22) : $signed(_GEN_26003); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26604 = 6'ha == state ? $signed(w_23) : $signed(_GEN_26004); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26605 = 6'ha == state ? $signed(w_24) : $signed(_GEN_26005); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26606 = 6'ha == state ? $signed(w_25) : $signed(_GEN_26006); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26607 = 6'ha == state ? $signed(w_26) : $signed(_GEN_26007); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26608 = 6'ha == state ? $signed(w_27) : $signed(_GEN_26008); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26609 = 6'ha == state ? $signed(w_28) : $signed(_GEN_26009); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26610 = 6'ha == state ? $signed(w_29) : $signed(_GEN_26010); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26611 = 6'ha == state ? $signed(w_30) : $signed(_GEN_26011); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26612 = 6'ha == state ? $signed(w_31) : $signed(_GEN_26012); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26613 = 6'ha == state ? $signed(w_32) : $signed(_GEN_26013); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26614 = 6'ha == state ? $signed(w_33) : $signed(_GEN_26014); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26615 = 6'ha == state ? $signed(w_34) : $signed(_GEN_26015); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26616 = 6'ha == state ? $signed(w_35) : $signed(_GEN_26016); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26617 = 6'ha == state ? $signed(w_36) : $signed(_GEN_26017); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26618 = 6'ha == state ? $signed(w_37) : $signed(_GEN_26018); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26619 = 6'ha == state ? $signed(w_38) : $signed(_GEN_26019); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26620 = 6'ha == state ? $signed(w_39) : $signed(_GEN_26020); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26621 = 6'ha == state ? $signed(w_40) : $signed(_GEN_26021); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26622 = 6'ha == state ? $signed(w_41) : $signed(_GEN_26022); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26623 = 6'ha == state ? $signed(w_42) : $signed(_GEN_26023); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26624 = 6'ha == state ? $signed(w_43) : $signed(_GEN_26024); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26625 = 6'ha == state ? $signed(w_44) : $signed(_GEN_26025); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26626 = 6'ha == state ? $signed(w_45) : $signed(_GEN_26026); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26627 = 6'ha == state ? $signed(w_46) : $signed(_GEN_26027); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26628 = 6'ha == state ? $signed(w_47) : $signed(_GEN_26028); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26629 = 6'ha == state ? $signed(w_48) : $signed(_GEN_26029); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26630 = 6'ha == state ? $signed(w_49) : $signed(_GEN_26030); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26631 = 6'ha == state ? $signed(w_50) : $signed(_GEN_26031); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26632 = 6'ha == state ? $signed(w_51) : $signed(_GEN_26032); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26633 = 6'ha == state ? $signed(w_52) : $signed(_GEN_26033); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26634 = 6'ha == state ? $signed(w_53) : $signed(_GEN_26034); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26635 = 6'ha == state ? $signed(w_54) : $signed(_GEN_26035); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26636 = 6'ha == state ? $signed(w_55) : $signed(_GEN_26036); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26637 = 6'ha == state ? $signed(w_56) : $signed(_GEN_26037); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26638 = 6'ha == state ? $signed(w_57) : $signed(_GEN_26038); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26639 = 6'ha == state ? $signed(w_58) : $signed(_GEN_26039); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26640 = 6'ha == state ? $signed(w_59) : $signed(_GEN_26040); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26641 = 6'ha == state ? $signed(w_60) : $signed(_GEN_26041); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26642 = 6'ha == state ? $signed(w_61) : $signed(_GEN_26042); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26643 = 6'ha == state ? $signed(w_62) : $signed(_GEN_26043); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26644 = 6'ha == state ? $signed(w_63) : $signed(_GEN_26044); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26645 = 6'ha == state ? $signed(w_64) : $signed(_GEN_26045); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26646 = 6'ha == state ? $signed(w_65) : $signed(_GEN_26046); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26647 = 6'ha == state ? $signed(w_66) : $signed(_GEN_26047); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26648 = 6'ha == state ? $signed(w_67) : $signed(_GEN_26048); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26649 = 6'ha == state ? $signed(w_68) : $signed(_GEN_26049); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26650 = 6'ha == state ? $signed(w_69) : $signed(_GEN_26050); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26651 = 6'ha == state ? $signed(w_70) : $signed(_GEN_26051); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26652 = 6'ha == state ? $signed(w_71) : $signed(_GEN_26052); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26653 = 6'ha == state ? $signed(w_72) : $signed(_GEN_26053); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26654 = 6'ha == state ? $signed(w_73) : $signed(_GEN_26054); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26655 = 6'ha == state ? $signed(w_74) : $signed(_GEN_26055); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26656 = 6'ha == state ? $signed(w_75) : $signed(_GEN_26056); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26657 = 6'ha == state ? $signed(w_76) : $signed(_GEN_26057); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26658 = 6'ha == state ? $signed(w_77) : $signed(_GEN_26058); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26659 = 6'ha == state ? $signed(w_78) : $signed(_GEN_26059); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26660 = 6'ha == state ? $signed(w_79) : $signed(_GEN_26060); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_26661 = 6'ha == state ? $signed(temp) : $signed(_GEN_26061); // @[digest.scala 38:19 81:19]
  wire  _GEN_26662 = 6'ha == state ? 1'h0 : _GEN_26062; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_26665 = 6'ha == state ? $signed(t) : $signed(_GEN_26065); // @[digest.scala 35:16 81:19]
  wire  _GEN_26666 = 6'ha == state ? 1'h0 : _GEN_26066; // @[digest.scala 81:19 48:24]
  wire  _GEN_26669 = 6'ha == state ? 1'h0 : _GEN_26069; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_26753 = 6'ha == state ? $signed(digest_0) : $signed(_GEN_26154); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26754 = 6'ha == state ? $signed(digest_1) : $signed(_GEN_26155); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26755 = 6'ha == state ? $signed(digest_2) : $signed(_GEN_26156); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26756 = 6'ha == state ? $signed(digest_3) : $signed(_GEN_26157); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26757 = 6'ha == state ? $signed(digest_4) : $signed(_GEN_26158); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26758 = 6'ha == state ? $signed(digest_5) : $signed(_GEN_26159); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26759 = 6'ha == state ? $signed(digest_6) : $signed(_GEN_26160); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26760 = 6'ha == state ? $signed(digest_7) : $signed(_GEN_26161); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26761 = 6'ha == state ? $signed(digest_8) : $signed(_GEN_26162); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26762 = 6'ha == state ? $signed(digest_9) : $signed(_GEN_26163); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26763 = 6'ha == state ? $signed(digest_10) : $signed(_GEN_26164); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26764 = 6'ha == state ? $signed(digest_11) : $signed(_GEN_26165); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26765 = 6'ha == state ? $signed(digest_12) : $signed(_GEN_26166); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26766 = 6'ha == state ? $signed(digest_13) : $signed(_GEN_26167); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26767 = 6'ha == state ? $signed(digest_14) : $signed(_GEN_26168); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26768 = 6'ha == state ? $signed(digest_15) : $signed(_GEN_26169); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26769 = 6'ha == state ? $signed(digest_16) : $signed(_GEN_26170); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26770 = 6'ha == state ? $signed(digest_17) : $signed(_GEN_26171); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26771 = 6'ha == state ? $signed(digest_18) : $signed(_GEN_26172); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26772 = 6'ha == state ? $signed(digest_19) : $signed(_GEN_26173); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26773 = 6'ha == state ? $signed(digest_20) : $signed(_GEN_26174); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26774 = 6'ha == state ? $signed(digest_21) : $signed(_GEN_26175); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26775 = 6'ha == state ? $signed(digest_22) : $signed(_GEN_26176); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26776 = 6'ha == state ? $signed(digest_23) : $signed(_GEN_26177); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26777 = 6'ha == state ? $signed(digest_24) : $signed(_GEN_26178); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26778 = 6'ha == state ? $signed(digest_25) : $signed(_GEN_26179); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26779 = 6'ha == state ? $signed(digest_26) : $signed(_GEN_26180); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26780 = 6'ha == state ? $signed(digest_27) : $signed(_GEN_26181); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26781 = 6'ha == state ? $signed(digest_28) : $signed(_GEN_26182); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26782 = 6'ha == state ? $signed(digest_29) : $signed(_GEN_26183); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26783 = 6'ha == state ? $signed(digest_30) : $signed(_GEN_26184); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26784 = 6'ha == state ? $signed(digest_31) : $signed(_GEN_26185); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26785 = 6'ha == state ? $signed(digest_32) : $signed(_GEN_26186); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26786 = 6'ha == state ? $signed(digest_33) : $signed(_GEN_26187); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26787 = 6'ha == state ? $signed(digest_34) : $signed(_GEN_26188); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26788 = 6'ha == state ? $signed(digest_35) : $signed(_GEN_26189); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26789 = 6'ha == state ? $signed(digest_36) : $signed(_GEN_26190); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26790 = 6'ha == state ? $signed(digest_37) : $signed(_GEN_26191); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26791 = 6'ha == state ? $signed(digest_38) : $signed(_GEN_26192); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26792 = 6'ha == state ? $signed(digest_39) : $signed(_GEN_26193); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26793 = 6'ha == state ? $signed(digest_40) : $signed(_GEN_26194); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26794 = 6'ha == state ? $signed(digest_41) : $signed(_GEN_26195); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26795 = 6'ha == state ? $signed(digest_42) : $signed(_GEN_26196); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26796 = 6'ha == state ? $signed(digest_43) : $signed(_GEN_26197); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26797 = 6'ha == state ? $signed(digest_44) : $signed(_GEN_26198); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26798 = 6'ha == state ? $signed(digest_45) : $signed(_GEN_26199); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26799 = 6'ha == state ? $signed(digest_46) : $signed(_GEN_26200); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26800 = 6'ha == state ? $signed(digest_47) : $signed(_GEN_26201); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26801 = 6'ha == state ? $signed(digest_48) : $signed(_GEN_26202); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26802 = 6'ha == state ? $signed(digest_49) : $signed(_GEN_26203); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26803 = 6'ha == state ? $signed(digest_50) : $signed(_GEN_26204); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26804 = 6'ha == state ? $signed(digest_51) : $signed(_GEN_26205); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26805 = 6'ha == state ? $signed(digest_52) : $signed(_GEN_26206); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26806 = 6'ha == state ? $signed(digest_53) : $signed(_GEN_26207); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26807 = 6'ha == state ? $signed(digest_54) : $signed(_GEN_26208); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26808 = 6'ha == state ? $signed(digest_55) : $signed(_GEN_26209); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26809 = 6'ha == state ? $signed(digest_56) : $signed(_GEN_26210); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26810 = 6'ha == state ? $signed(digest_57) : $signed(_GEN_26211); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26811 = 6'ha == state ? $signed(digest_58) : $signed(_GEN_26212); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26812 = 6'ha == state ? $signed(digest_59) : $signed(_GEN_26213); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26813 = 6'ha == state ? $signed(digest_60) : $signed(_GEN_26214); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26814 = 6'ha == state ? $signed(digest_61) : $signed(_GEN_26215); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26815 = 6'ha == state ? $signed(digest_62) : $signed(_GEN_26216); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26816 = 6'ha == state ? $signed(digest_63) : $signed(_GEN_26217); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26817 = 6'ha == state ? $signed(digest_64) : $signed(_GEN_26218); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26818 = 6'ha == state ? $signed(digest_65) : $signed(_GEN_26219); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26819 = 6'ha == state ? $signed(digest_66) : $signed(_GEN_26220); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26820 = 6'ha == state ? $signed(digest_67) : $signed(_GEN_26221); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26821 = 6'ha == state ? $signed(digest_68) : $signed(_GEN_26222); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26822 = 6'ha == state ? $signed(digest_69) : $signed(_GEN_26223); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26823 = 6'ha == state ? $signed(digest_70) : $signed(_GEN_26224); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26824 = 6'ha == state ? $signed(digest_71) : $signed(_GEN_26225); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26825 = 6'ha == state ? $signed(digest_72) : $signed(_GEN_26226); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26826 = 6'ha == state ? $signed(digest_73) : $signed(_GEN_26227); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26827 = 6'ha == state ? $signed(digest_74) : $signed(_GEN_26228); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26828 = 6'ha == state ? $signed(digest_75) : $signed(_GEN_26229); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26829 = 6'ha == state ? $signed(digest_76) : $signed(_GEN_26230); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26830 = 6'ha == state ? $signed(digest_77) : $signed(_GEN_26231); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26831 = 6'ha == state ? $signed(digest_78) : $signed(_GEN_26232); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_26832 = 6'ha == state ? $signed(digest_79) : $signed(_GEN_26233); // @[digest.scala 81:19 53:21]
  wire  _GEN_26834 = 6'ha == state ? 1'h0 : _GEN_26235; // @[digest.scala 81:19 58:25]
  wire  _GEN_26917 = 6'ha == state ? 1'h0 : _GEN_26318; // @[digest.scala 81:19 63:25]
  wire  _GEN_27000 = 6'ha == state ? 1'h0 : _GEN_26401; // @[digest.scala 81:19 68:25]
  wire  _GEN_27083 = 6'ha == state ? 1'h0 : _GEN_26484; // @[digest.scala 81:19 73:25]
  wire  _GEN_27166 = 6'ha == state ? 1'h0 : _GEN_26567; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_27167 = 6'h9 == state ? $signed(_GEN_481) : $signed(blks_0); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27168 = 6'h9 == state ? $signed(_GEN_482) : $signed(blks_1); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27169 = 6'h9 == state ? $signed(_GEN_483) : $signed(blks_2); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27170 = 6'h9 == state ? $signed(_GEN_484) : $signed(blks_3); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27171 = 6'h9 == state ? $signed(_GEN_485) : $signed(blks_4); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27172 = 6'h9 == state ? $signed(_GEN_486) : $signed(blks_5); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27173 = 6'h9 == state ? $signed(_GEN_487) : $signed(blks_6); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27174 = 6'h9 == state ? $signed(_GEN_488) : $signed(blks_7); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27175 = 6'h9 == state ? $signed(_GEN_489) : $signed(blks_8); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27176 = 6'h9 == state ? $signed(_GEN_490) : $signed(blks_9); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27177 = 6'h9 == state ? $signed(_GEN_491) : $signed(blks_10); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27178 = 6'h9 == state ? $signed(_GEN_492) : $signed(blks_11); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27179 = 6'h9 == state ? $signed(_GEN_493) : $signed(blks_12); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27180 = 6'h9 == state ? $signed(_GEN_494) : $signed(blks_13); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27181 = 6'h9 == state ? $signed(_GEN_495) : $signed(blks_14); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27182 = 6'h9 == state ? $signed(_GEN_496) : $signed(blks_15); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27183 = 6'h9 == state ? $signed(_GEN_497) : $signed(blks_16); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27184 = 6'h9 == state ? $signed(_GEN_498) : $signed(blks_17); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27185 = 6'h9 == state ? $signed(_GEN_499) : $signed(blks_18); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27186 = 6'h9 == state ? $signed(_GEN_500) : $signed(blks_19); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27187 = 6'h9 == state ? $signed(_GEN_501) : $signed(blks_20); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27188 = 6'h9 == state ? $signed(_GEN_502) : $signed(blks_21); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27189 = 6'h9 == state ? $signed(_GEN_503) : $signed(blks_22); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27190 = 6'h9 == state ? $signed(_GEN_504) : $signed(blks_23); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27191 = 6'h9 == state ? $signed(_GEN_505) : $signed(blks_24); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27192 = 6'h9 == state ? $signed(_GEN_506) : $signed(blks_25); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27193 = 6'h9 == state ? $signed(_GEN_507) : $signed(blks_26); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27194 = 6'h9 == state ? $signed(_GEN_508) : $signed(blks_27); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27195 = 6'h9 == state ? $signed(_GEN_509) : $signed(blks_28); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27196 = 6'h9 == state ? $signed(_GEN_510) : $signed(blks_29); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27197 = 6'h9 == state ? $signed(_GEN_511) : $signed(blks_30); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27198 = 6'h9 == state ? $signed(_GEN_512) : $signed(blks_31); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27199 = 6'h9 == state ? $signed(_GEN_513) : $signed(blks_32); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27200 = 6'h9 == state ? $signed(_GEN_514) : $signed(blks_33); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27201 = 6'h9 == state ? $signed(_GEN_515) : $signed(blks_34); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27202 = 6'h9 == state ? $signed(_GEN_516) : $signed(blks_35); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27203 = 6'h9 == state ? $signed(_GEN_517) : $signed(blks_36); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27204 = 6'h9 == state ? $signed(_GEN_518) : $signed(blks_37); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27205 = 6'h9 == state ? $signed(_GEN_519) : $signed(blks_38); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27206 = 6'h9 == state ? $signed(_GEN_520) : $signed(blks_39); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27207 = 6'h9 == state ? $signed(_GEN_521) : $signed(blks_40); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27208 = 6'h9 == state ? $signed(_GEN_522) : $signed(blks_41); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27209 = 6'h9 == state ? $signed(_GEN_523) : $signed(blks_42); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27210 = 6'h9 == state ? $signed(_GEN_524) : $signed(blks_43); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27211 = 6'h9 == state ? $signed(_GEN_525) : $signed(blks_44); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27212 = 6'h9 == state ? $signed(_GEN_526) : $signed(blks_45); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27213 = 6'h9 == state ? $signed(_GEN_527) : $signed(blks_46); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27214 = 6'h9 == state ? $signed(_GEN_528) : $signed(blks_47); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27215 = 6'h9 == state ? $signed(_GEN_529) : $signed(blks_48); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27216 = 6'h9 == state ? $signed(_GEN_530) : $signed(blks_49); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27217 = 6'h9 == state ? $signed(_GEN_531) : $signed(blks_50); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27218 = 6'h9 == state ? $signed(_GEN_532) : $signed(blks_51); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27219 = 6'h9 == state ? $signed(_GEN_533) : $signed(blks_52); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27220 = 6'h9 == state ? $signed(_GEN_534) : $signed(blks_53); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27221 = 6'h9 == state ? $signed(_GEN_535) : $signed(blks_54); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27222 = 6'h9 == state ? $signed(_GEN_536) : $signed(blks_55); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27223 = 6'h9 == state ? $signed(_GEN_537) : $signed(blks_56); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27224 = 6'h9 == state ? $signed(_GEN_538) : $signed(blks_57); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27225 = 6'h9 == state ? $signed(_GEN_539) : $signed(blks_58); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27226 = 6'h9 == state ? $signed(_GEN_540) : $signed(blks_59); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27227 = 6'h9 == state ? $signed(_GEN_541) : $signed(blks_60); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27228 = 6'h9 == state ? $signed(_GEN_542) : $signed(blks_61); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27229 = 6'h9 == state ? $signed(_GEN_543) : $signed(blks_62); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27230 = 6'h9 == state ? $signed(_GEN_544) : $signed(blks_63); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27231 = 6'h9 == state ? $signed(_GEN_545) : $signed(blks_64); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27232 = 6'h9 == state ? $signed(_GEN_546) : $signed(blks_65); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27233 = 6'h9 == state ? $signed(_GEN_547) : $signed(blks_66); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27234 = 6'h9 == state ? $signed(_GEN_548) : $signed(blks_67); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27235 = 6'h9 == state ? $signed(_GEN_549) : $signed(blks_68); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27236 = 6'h9 == state ? $signed(_GEN_550) : $signed(blks_69); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27237 = 6'h9 == state ? $signed(_GEN_551) : $signed(blks_70); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27238 = 6'h9 == state ? $signed(_GEN_552) : $signed(blks_71); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27239 = 6'h9 == state ? $signed(_GEN_553) : $signed(blks_72); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27240 = 6'h9 == state ? $signed(_GEN_554) : $signed(blks_73); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27241 = 6'h9 == state ? $signed(_GEN_555) : $signed(blks_74); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27242 = 6'h9 == state ? $signed(_GEN_556) : $signed(blks_75); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27243 = 6'h9 == state ? $signed(_GEN_557) : $signed(blks_76); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27244 = 6'h9 == state ? $signed(_GEN_558) : $signed(blks_77); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27245 = 6'h9 == state ? $signed(_GEN_559) : $signed(blks_78); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_27246 = 6'h9 == state ? $signed(_GEN_560) : $signed(blks_79); // @[digest.scala 39:19 81:19]
  wire [5:0] _GEN_27247 = 6'h9 == state ? 6'ha : _GEN_26569; // @[digest.scala 122:19 81:19]
  wire [31:0] _GEN_27248 = 6'h9 == state ? $signed(a) : $signed(_GEN_26568); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_27249 = 6'h9 == state ? $signed(b) : $signed(_GEN_26570); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_27250 = 6'h9 == state ? $signed(c) : $signed(_GEN_26571); // @[digest.scala 26:16 81:19]
  wire [31:0] _GEN_27251 = 6'h9 == state ? $signed(d) : $signed(_GEN_26572); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_27252 = 6'h9 == state ? $signed(e) : $signed(_GEN_26573); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_27253 = 6'h9 == state ? $signed(i) : $signed(_GEN_26574); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_27254 = 6'h9 == state ? $signed(olda) : $signed(_GEN_26575); // @[digest.scala 29:19 81:19]
  wire [31:0] _GEN_27255 = 6'h9 == state ? $signed(oldb) : $signed(_GEN_26576); // @[digest.scala 30:19 81:19]
  wire [31:0] _GEN_27256 = 6'h9 == state ? $signed(oldc) : $signed(_GEN_26577); // @[digest.scala 31:19 81:19]
  wire [31:0] _GEN_27257 = 6'h9 == state ? $signed(oldd) : $signed(_GEN_26578); // @[digest.scala 32:19 81:19]
  wire [31:0] _GEN_27258 = 6'h9 == state ? $signed(olde) : $signed(_GEN_26579); // @[digest.scala 33:19 81:19]
  wire [31:0] _GEN_27259 = 6'h9 == state ? $signed(j) : $signed(_GEN_26580); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_27260 = 6'h9 == state ? $signed(w_0) : $signed(_GEN_26581); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27261 = 6'h9 == state ? $signed(w_1) : $signed(_GEN_26582); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27262 = 6'h9 == state ? $signed(w_2) : $signed(_GEN_26583); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27263 = 6'h9 == state ? $signed(w_3) : $signed(_GEN_26584); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27264 = 6'h9 == state ? $signed(w_4) : $signed(_GEN_26585); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27265 = 6'h9 == state ? $signed(w_5) : $signed(_GEN_26586); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27266 = 6'h9 == state ? $signed(w_6) : $signed(_GEN_26587); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27267 = 6'h9 == state ? $signed(w_7) : $signed(_GEN_26588); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27268 = 6'h9 == state ? $signed(w_8) : $signed(_GEN_26589); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27269 = 6'h9 == state ? $signed(w_9) : $signed(_GEN_26590); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27270 = 6'h9 == state ? $signed(w_10) : $signed(_GEN_26591); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27271 = 6'h9 == state ? $signed(w_11) : $signed(_GEN_26592); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27272 = 6'h9 == state ? $signed(w_12) : $signed(_GEN_26593); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27273 = 6'h9 == state ? $signed(w_13) : $signed(_GEN_26594); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27274 = 6'h9 == state ? $signed(w_14) : $signed(_GEN_26595); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27275 = 6'h9 == state ? $signed(w_15) : $signed(_GEN_26596); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27276 = 6'h9 == state ? $signed(w_16) : $signed(_GEN_26597); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27277 = 6'h9 == state ? $signed(w_17) : $signed(_GEN_26598); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27278 = 6'h9 == state ? $signed(w_18) : $signed(_GEN_26599); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27279 = 6'h9 == state ? $signed(w_19) : $signed(_GEN_26600); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27280 = 6'h9 == state ? $signed(w_20) : $signed(_GEN_26601); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27281 = 6'h9 == state ? $signed(w_21) : $signed(_GEN_26602); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27282 = 6'h9 == state ? $signed(w_22) : $signed(_GEN_26603); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27283 = 6'h9 == state ? $signed(w_23) : $signed(_GEN_26604); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27284 = 6'h9 == state ? $signed(w_24) : $signed(_GEN_26605); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27285 = 6'h9 == state ? $signed(w_25) : $signed(_GEN_26606); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27286 = 6'h9 == state ? $signed(w_26) : $signed(_GEN_26607); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27287 = 6'h9 == state ? $signed(w_27) : $signed(_GEN_26608); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27288 = 6'h9 == state ? $signed(w_28) : $signed(_GEN_26609); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27289 = 6'h9 == state ? $signed(w_29) : $signed(_GEN_26610); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27290 = 6'h9 == state ? $signed(w_30) : $signed(_GEN_26611); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27291 = 6'h9 == state ? $signed(w_31) : $signed(_GEN_26612); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27292 = 6'h9 == state ? $signed(w_32) : $signed(_GEN_26613); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27293 = 6'h9 == state ? $signed(w_33) : $signed(_GEN_26614); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27294 = 6'h9 == state ? $signed(w_34) : $signed(_GEN_26615); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27295 = 6'h9 == state ? $signed(w_35) : $signed(_GEN_26616); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27296 = 6'h9 == state ? $signed(w_36) : $signed(_GEN_26617); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27297 = 6'h9 == state ? $signed(w_37) : $signed(_GEN_26618); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27298 = 6'h9 == state ? $signed(w_38) : $signed(_GEN_26619); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27299 = 6'h9 == state ? $signed(w_39) : $signed(_GEN_26620); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27300 = 6'h9 == state ? $signed(w_40) : $signed(_GEN_26621); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27301 = 6'h9 == state ? $signed(w_41) : $signed(_GEN_26622); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27302 = 6'h9 == state ? $signed(w_42) : $signed(_GEN_26623); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27303 = 6'h9 == state ? $signed(w_43) : $signed(_GEN_26624); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27304 = 6'h9 == state ? $signed(w_44) : $signed(_GEN_26625); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27305 = 6'h9 == state ? $signed(w_45) : $signed(_GEN_26626); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27306 = 6'h9 == state ? $signed(w_46) : $signed(_GEN_26627); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27307 = 6'h9 == state ? $signed(w_47) : $signed(_GEN_26628); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27308 = 6'h9 == state ? $signed(w_48) : $signed(_GEN_26629); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27309 = 6'h9 == state ? $signed(w_49) : $signed(_GEN_26630); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27310 = 6'h9 == state ? $signed(w_50) : $signed(_GEN_26631); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27311 = 6'h9 == state ? $signed(w_51) : $signed(_GEN_26632); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27312 = 6'h9 == state ? $signed(w_52) : $signed(_GEN_26633); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27313 = 6'h9 == state ? $signed(w_53) : $signed(_GEN_26634); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27314 = 6'h9 == state ? $signed(w_54) : $signed(_GEN_26635); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27315 = 6'h9 == state ? $signed(w_55) : $signed(_GEN_26636); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27316 = 6'h9 == state ? $signed(w_56) : $signed(_GEN_26637); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27317 = 6'h9 == state ? $signed(w_57) : $signed(_GEN_26638); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27318 = 6'h9 == state ? $signed(w_58) : $signed(_GEN_26639); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27319 = 6'h9 == state ? $signed(w_59) : $signed(_GEN_26640); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27320 = 6'h9 == state ? $signed(w_60) : $signed(_GEN_26641); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27321 = 6'h9 == state ? $signed(w_61) : $signed(_GEN_26642); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27322 = 6'h9 == state ? $signed(w_62) : $signed(_GEN_26643); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27323 = 6'h9 == state ? $signed(w_63) : $signed(_GEN_26644); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27324 = 6'h9 == state ? $signed(w_64) : $signed(_GEN_26645); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27325 = 6'h9 == state ? $signed(w_65) : $signed(_GEN_26646); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27326 = 6'h9 == state ? $signed(w_66) : $signed(_GEN_26647); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27327 = 6'h9 == state ? $signed(w_67) : $signed(_GEN_26648); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27328 = 6'h9 == state ? $signed(w_68) : $signed(_GEN_26649); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27329 = 6'h9 == state ? $signed(w_69) : $signed(_GEN_26650); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27330 = 6'h9 == state ? $signed(w_70) : $signed(_GEN_26651); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27331 = 6'h9 == state ? $signed(w_71) : $signed(_GEN_26652); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27332 = 6'h9 == state ? $signed(w_72) : $signed(_GEN_26653); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27333 = 6'h9 == state ? $signed(w_73) : $signed(_GEN_26654); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27334 = 6'h9 == state ? $signed(w_74) : $signed(_GEN_26655); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27335 = 6'h9 == state ? $signed(w_75) : $signed(_GEN_26656); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27336 = 6'h9 == state ? $signed(w_76) : $signed(_GEN_26657); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27337 = 6'h9 == state ? $signed(w_77) : $signed(_GEN_26658); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27338 = 6'h9 == state ? $signed(w_78) : $signed(_GEN_26659); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27339 = 6'h9 == state ? $signed(w_79) : $signed(_GEN_26660); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27340 = 6'h9 == state ? $signed(temp) : $signed(_GEN_26661); // @[digest.scala 38:19 81:19]
  wire  _GEN_27341 = 6'h9 == state ? 1'h0 : _GEN_26662; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_27344 = 6'h9 == state ? $signed(t) : $signed(_GEN_26665); // @[digest.scala 35:16 81:19]
  wire  _GEN_27345 = 6'h9 == state ? 1'h0 : _GEN_26666; // @[digest.scala 81:19 48:24]
  wire  _GEN_27348 = 6'h9 == state ? 1'h0 : _GEN_26669; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_27432 = 6'h9 == state ? $signed(digest_0) : $signed(_GEN_26753); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27433 = 6'h9 == state ? $signed(digest_1) : $signed(_GEN_26754); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27434 = 6'h9 == state ? $signed(digest_2) : $signed(_GEN_26755); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27435 = 6'h9 == state ? $signed(digest_3) : $signed(_GEN_26756); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27436 = 6'h9 == state ? $signed(digest_4) : $signed(_GEN_26757); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27437 = 6'h9 == state ? $signed(digest_5) : $signed(_GEN_26758); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27438 = 6'h9 == state ? $signed(digest_6) : $signed(_GEN_26759); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27439 = 6'h9 == state ? $signed(digest_7) : $signed(_GEN_26760); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27440 = 6'h9 == state ? $signed(digest_8) : $signed(_GEN_26761); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27441 = 6'h9 == state ? $signed(digest_9) : $signed(_GEN_26762); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27442 = 6'h9 == state ? $signed(digest_10) : $signed(_GEN_26763); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27443 = 6'h9 == state ? $signed(digest_11) : $signed(_GEN_26764); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27444 = 6'h9 == state ? $signed(digest_12) : $signed(_GEN_26765); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27445 = 6'h9 == state ? $signed(digest_13) : $signed(_GEN_26766); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27446 = 6'h9 == state ? $signed(digest_14) : $signed(_GEN_26767); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27447 = 6'h9 == state ? $signed(digest_15) : $signed(_GEN_26768); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27448 = 6'h9 == state ? $signed(digest_16) : $signed(_GEN_26769); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27449 = 6'h9 == state ? $signed(digest_17) : $signed(_GEN_26770); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27450 = 6'h9 == state ? $signed(digest_18) : $signed(_GEN_26771); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27451 = 6'h9 == state ? $signed(digest_19) : $signed(_GEN_26772); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27452 = 6'h9 == state ? $signed(digest_20) : $signed(_GEN_26773); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27453 = 6'h9 == state ? $signed(digest_21) : $signed(_GEN_26774); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27454 = 6'h9 == state ? $signed(digest_22) : $signed(_GEN_26775); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27455 = 6'h9 == state ? $signed(digest_23) : $signed(_GEN_26776); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27456 = 6'h9 == state ? $signed(digest_24) : $signed(_GEN_26777); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27457 = 6'h9 == state ? $signed(digest_25) : $signed(_GEN_26778); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27458 = 6'h9 == state ? $signed(digest_26) : $signed(_GEN_26779); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27459 = 6'h9 == state ? $signed(digest_27) : $signed(_GEN_26780); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27460 = 6'h9 == state ? $signed(digest_28) : $signed(_GEN_26781); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27461 = 6'h9 == state ? $signed(digest_29) : $signed(_GEN_26782); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27462 = 6'h9 == state ? $signed(digest_30) : $signed(_GEN_26783); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27463 = 6'h9 == state ? $signed(digest_31) : $signed(_GEN_26784); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27464 = 6'h9 == state ? $signed(digest_32) : $signed(_GEN_26785); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27465 = 6'h9 == state ? $signed(digest_33) : $signed(_GEN_26786); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27466 = 6'h9 == state ? $signed(digest_34) : $signed(_GEN_26787); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27467 = 6'h9 == state ? $signed(digest_35) : $signed(_GEN_26788); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27468 = 6'h9 == state ? $signed(digest_36) : $signed(_GEN_26789); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27469 = 6'h9 == state ? $signed(digest_37) : $signed(_GEN_26790); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27470 = 6'h9 == state ? $signed(digest_38) : $signed(_GEN_26791); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27471 = 6'h9 == state ? $signed(digest_39) : $signed(_GEN_26792); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27472 = 6'h9 == state ? $signed(digest_40) : $signed(_GEN_26793); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27473 = 6'h9 == state ? $signed(digest_41) : $signed(_GEN_26794); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27474 = 6'h9 == state ? $signed(digest_42) : $signed(_GEN_26795); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27475 = 6'h9 == state ? $signed(digest_43) : $signed(_GEN_26796); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27476 = 6'h9 == state ? $signed(digest_44) : $signed(_GEN_26797); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27477 = 6'h9 == state ? $signed(digest_45) : $signed(_GEN_26798); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27478 = 6'h9 == state ? $signed(digest_46) : $signed(_GEN_26799); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27479 = 6'h9 == state ? $signed(digest_47) : $signed(_GEN_26800); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27480 = 6'h9 == state ? $signed(digest_48) : $signed(_GEN_26801); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27481 = 6'h9 == state ? $signed(digest_49) : $signed(_GEN_26802); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27482 = 6'h9 == state ? $signed(digest_50) : $signed(_GEN_26803); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27483 = 6'h9 == state ? $signed(digest_51) : $signed(_GEN_26804); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27484 = 6'h9 == state ? $signed(digest_52) : $signed(_GEN_26805); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27485 = 6'h9 == state ? $signed(digest_53) : $signed(_GEN_26806); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27486 = 6'h9 == state ? $signed(digest_54) : $signed(_GEN_26807); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27487 = 6'h9 == state ? $signed(digest_55) : $signed(_GEN_26808); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27488 = 6'h9 == state ? $signed(digest_56) : $signed(_GEN_26809); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27489 = 6'h9 == state ? $signed(digest_57) : $signed(_GEN_26810); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27490 = 6'h9 == state ? $signed(digest_58) : $signed(_GEN_26811); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27491 = 6'h9 == state ? $signed(digest_59) : $signed(_GEN_26812); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27492 = 6'h9 == state ? $signed(digest_60) : $signed(_GEN_26813); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27493 = 6'h9 == state ? $signed(digest_61) : $signed(_GEN_26814); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27494 = 6'h9 == state ? $signed(digest_62) : $signed(_GEN_26815); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27495 = 6'h9 == state ? $signed(digest_63) : $signed(_GEN_26816); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27496 = 6'h9 == state ? $signed(digest_64) : $signed(_GEN_26817); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27497 = 6'h9 == state ? $signed(digest_65) : $signed(_GEN_26818); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27498 = 6'h9 == state ? $signed(digest_66) : $signed(_GEN_26819); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27499 = 6'h9 == state ? $signed(digest_67) : $signed(_GEN_26820); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27500 = 6'h9 == state ? $signed(digest_68) : $signed(_GEN_26821); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27501 = 6'h9 == state ? $signed(digest_69) : $signed(_GEN_26822); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27502 = 6'h9 == state ? $signed(digest_70) : $signed(_GEN_26823); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27503 = 6'h9 == state ? $signed(digest_71) : $signed(_GEN_26824); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27504 = 6'h9 == state ? $signed(digest_72) : $signed(_GEN_26825); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27505 = 6'h9 == state ? $signed(digest_73) : $signed(_GEN_26826); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27506 = 6'h9 == state ? $signed(digest_74) : $signed(_GEN_26827); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27507 = 6'h9 == state ? $signed(digest_75) : $signed(_GEN_26828); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27508 = 6'h9 == state ? $signed(digest_76) : $signed(_GEN_26829); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27509 = 6'h9 == state ? $signed(digest_77) : $signed(_GEN_26830); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27510 = 6'h9 == state ? $signed(digest_78) : $signed(_GEN_26831); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_27511 = 6'h9 == state ? $signed(digest_79) : $signed(_GEN_26832); // @[digest.scala 81:19 53:21]
  wire  _GEN_27513 = 6'h9 == state ? 1'h0 : _GEN_26834; // @[digest.scala 81:19 58:25]
  wire  _GEN_27596 = 6'h9 == state ? 1'h0 : _GEN_26917; // @[digest.scala 81:19 63:25]
  wire  _GEN_27679 = 6'h9 == state ? 1'h0 : _GEN_27000; // @[digest.scala 81:19 68:25]
  wire  _GEN_27762 = 6'h9 == state ? 1'h0 : _GEN_27083; // @[digest.scala 81:19 73:25]
  wire  _GEN_27845 = 6'h9 == state ? 1'h0 : _GEN_27166; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_27846 = 6'h8 == state ? $signed(_GEN_241) : $signed(_GEN_27167); // @[digest.scala 81:19]
  wire [31:0] _GEN_27847 = 6'h8 == state ? $signed(_GEN_242) : $signed(_GEN_27168); // @[digest.scala 81:19]
  wire [31:0] _GEN_27848 = 6'h8 == state ? $signed(_GEN_243) : $signed(_GEN_27169); // @[digest.scala 81:19]
  wire [31:0] _GEN_27849 = 6'h8 == state ? $signed(_GEN_244) : $signed(_GEN_27170); // @[digest.scala 81:19]
  wire [31:0] _GEN_27850 = 6'h8 == state ? $signed(_GEN_245) : $signed(_GEN_27171); // @[digest.scala 81:19]
  wire [31:0] _GEN_27851 = 6'h8 == state ? $signed(_GEN_246) : $signed(_GEN_27172); // @[digest.scala 81:19]
  wire [31:0] _GEN_27852 = 6'h8 == state ? $signed(_GEN_247) : $signed(_GEN_27173); // @[digest.scala 81:19]
  wire [31:0] _GEN_27853 = 6'h8 == state ? $signed(_GEN_248) : $signed(_GEN_27174); // @[digest.scala 81:19]
  wire [31:0] _GEN_27854 = 6'h8 == state ? $signed(_GEN_249) : $signed(_GEN_27175); // @[digest.scala 81:19]
  wire [31:0] _GEN_27855 = 6'h8 == state ? $signed(_GEN_250) : $signed(_GEN_27176); // @[digest.scala 81:19]
  wire [31:0] _GEN_27856 = 6'h8 == state ? $signed(_GEN_251) : $signed(_GEN_27177); // @[digest.scala 81:19]
  wire [31:0] _GEN_27857 = 6'h8 == state ? $signed(_GEN_252) : $signed(_GEN_27178); // @[digest.scala 81:19]
  wire [31:0] _GEN_27858 = 6'h8 == state ? $signed(_GEN_253) : $signed(_GEN_27179); // @[digest.scala 81:19]
  wire [31:0] _GEN_27859 = 6'h8 == state ? $signed(_GEN_254) : $signed(_GEN_27180); // @[digest.scala 81:19]
  wire [31:0] _GEN_27860 = 6'h8 == state ? $signed(_GEN_255) : $signed(_GEN_27181); // @[digest.scala 81:19]
  wire [31:0] _GEN_27861 = 6'h8 == state ? $signed(_GEN_256) : $signed(_GEN_27182); // @[digest.scala 81:19]
  wire [31:0] _GEN_27862 = 6'h8 == state ? $signed(_GEN_257) : $signed(_GEN_27183); // @[digest.scala 81:19]
  wire [31:0] _GEN_27863 = 6'h8 == state ? $signed(_GEN_258) : $signed(_GEN_27184); // @[digest.scala 81:19]
  wire [31:0] _GEN_27864 = 6'h8 == state ? $signed(_GEN_259) : $signed(_GEN_27185); // @[digest.scala 81:19]
  wire [31:0] _GEN_27865 = 6'h8 == state ? $signed(_GEN_260) : $signed(_GEN_27186); // @[digest.scala 81:19]
  wire [31:0] _GEN_27866 = 6'h8 == state ? $signed(_GEN_261) : $signed(_GEN_27187); // @[digest.scala 81:19]
  wire [31:0] _GEN_27867 = 6'h8 == state ? $signed(_GEN_262) : $signed(_GEN_27188); // @[digest.scala 81:19]
  wire [31:0] _GEN_27868 = 6'h8 == state ? $signed(_GEN_263) : $signed(_GEN_27189); // @[digest.scala 81:19]
  wire [31:0] _GEN_27869 = 6'h8 == state ? $signed(_GEN_264) : $signed(_GEN_27190); // @[digest.scala 81:19]
  wire [31:0] _GEN_27870 = 6'h8 == state ? $signed(_GEN_265) : $signed(_GEN_27191); // @[digest.scala 81:19]
  wire [31:0] _GEN_27871 = 6'h8 == state ? $signed(_GEN_266) : $signed(_GEN_27192); // @[digest.scala 81:19]
  wire [31:0] _GEN_27872 = 6'h8 == state ? $signed(_GEN_267) : $signed(_GEN_27193); // @[digest.scala 81:19]
  wire [31:0] _GEN_27873 = 6'h8 == state ? $signed(_GEN_268) : $signed(_GEN_27194); // @[digest.scala 81:19]
  wire [31:0] _GEN_27874 = 6'h8 == state ? $signed(_GEN_269) : $signed(_GEN_27195); // @[digest.scala 81:19]
  wire [31:0] _GEN_27875 = 6'h8 == state ? $signed(_GEN_270) : $signed(_GEN_27196); // @[digest.scala 81:19]
  wire [31:0] _GEN_27876 = 6'h8 == state ? $signed(_GEN_271) : $signed(_GEN_27197); // @[digest.scala 81:19]
  wire [31:0] _GEN_27877 = 6'h8 == state ? $signed(_GEN_272) : $signed(_GEN_27198); // @[digest.scala 81:19]
  wire [31:0] _GEN_27878 = 6'h8 == state ? $signed(_GEN_273) : $signed(_GEN_27199); // @[digest.scala 81:19]
  wire [31:0] _GEN_27879 = 6'h8 == state ? $signed(_GEN_274) : $signed(_GEN_27200); // @[digest.scala 81:19]
  wire [31:0] _GEN_27880 = 6'h8 == state ? $signed(_GEN_275) : $signed(_GEN_27201); // @[digest.scala 81:19]
  wire [31:0] _GEN_27881 = 6'h8 == state ? $signed(_GEN_276) : $signed(_GEN_27202); // @[digest.scala 81:19]
  wire [31:0] _GEN_27882 = 6'h8 == state ? $signed(_GEN_277) : $signed(_GEN_27203); // @[digest.scala 81:19]
  wire [31:0] _GEN_27883 = 6'h8 == state ? $signed(_GEN_278) : $signed(_GEN_27204); // @[digest.scala 81:19]
  wire [31:0] _GEN_27884 = 6'h8 == state ? $signed(_GEN_279) : $signed(_GEN_27205); // @[digest.scala 81:19]
  wire [31:0] _GEN_27885 = 6'h8 == state ? $signed(_GEN_280) : $signed(_GEN_27206); // @[digest.scala 81:19]
  wire [31:0] _GEN_27886 = 6'h8 == state ? $signed(_GEN_281) : $signed(_GEN_27207); // @[digest.scala 81:19]
  wire [31:0] _GEN_27887 = 6'h8 == state ? $signed(_GEN_282) : $signed(_GEN_27208); // @[digest.scala 81:19]
  wire [31:0] _GEN_27888 = 6'h8 == state ? $signed(_GEN_283) : $signed(_GEN_27209); // @[digest.scala 81:19]
  wire [31:0] _GEN_27889 = 6'h8 == state ? $signed(_GEN_284) : $signed(_GEN_27210); // @[digest.scala 81:19]
  wire [31:0] _GEN_27890 = 6'h8 == state ? $signed(_GEN_285) : $signed(_GEN_27211); // @[digest.scala 81:19]
  wire [31:0] _GEN_27891 = 6'h8 == state ? $signed(_GEN_286) : $signed(_GEN_27212); // @[digest.scala 81:19]
  wire [31:0] _GEN_27892 = 6'h8 == state ? $signed(_GEN_287) : $signed(_GEN_27213); // @[digest.scala 81:19]
  wire [31:0] _GEN_27893 = 6'h8 == state ? $signed(_GEN_288) : $signed(_GEN_27214); // @[digest.scala 81:19]
  wire [31:0] _GEN_27894 = 6'h8 == state ? $signed(_GEN_289) : $signed(_GEN_27215); // @[digest.scala 81:19]
  wire [31:0] _GEN_27895 = 6'h8 == state ? $signed(_GEN_290) : $signed(_GEN_27216); // @[digest.scala 81:19]
  wire [31:0] _GEN_27896 = 6'h8 == state ? $signed(_GEN_291) : $signed(_GEN_27217); // @[digest.scala 81:19]
  wire [31:0] _GEN_27897 = 6'h8 == state ? $signed(_GEN_292) : $signed(_GEN_27218); // @[digest.scala 81:19]
  wire [31:0] _GEN_27898 = 6'h8 == state ? $signed(_GEN_293) : $signed(_GEN_27219); // @[digest.scala 81:19]
  wire [31:0] _GEN_27899 = 6'h8 == state ? $signed(_GEN_294) : $signed(_GEN_27220); // @[digest.scala 81:19]
  wire [31:0] _GEN_27900 = 6'h8 == state ? $signed(_GEN_295) : $signed(_GEN_27221); // @[digest.scala 81:19]
  wire [31:0] _GEN_27901 = 6'h8 == state ? $signed(_GEN_296) : $signed(_GEN_27222); // @[digest.scala 81:19]
  wire [31:0] _GEN_27902 = 6'h8 == state ? $signed(_GEN_297) : $signed(_GEN_27223); // @[digest.scala 81:19]
  wire [31:0] _GEN_27903 = 6'h8 == state ? $signed(_GEN_298) : $signed(_GEN_27224); // @[digest.scala 81:19]
  wire [31:0] _GEN_27904 = 6'h8 == state ? $signed(_GEN_299) : $signed(_GEN_27225); // @[digest.scala 81:19]
  wire [31:0] _GEN_27905 = 6'h8 == state ? $signed(_GEN_300) : $signed(_GEN_27226); // @[digest.scala 81:19]
  wire [31:0] _GEN_27906 = 6'h8 == state ? $signed(_GEN_301) : $signed(_GEN_27227); // @[digest.scala 81:19]
  wire [31:0] _GEN_27907 = 6'h8 == state ? $signed(_GEN_302) : $signed(_GEN_27228); // @[digest.scala 81:19]
  wire [31:0] _GEN_27908 = 6'h8 == state ? $signed(_GEN_303) : $signed(_GEN_27229); // @[digest.scala 81:19]
  wire [31:0] _GEN_27909 = 6'h8 == state ? $signed(_GEN_304) : $signed(_GEN_27230); // @[digest.scala 81:19]
  wire [31:0] _GEN_27910 = 6'h8 == state ? $signed(_GEN_305) : $signed(_GEN_27231); // @[digest.scala 81:19]
  wire [31:0] _GEN_27911 = 6'h8 == state ? $signed(_GEN_306) : $signed(_GEN_27232); // @[digest.scala 81:19]
  wire [31:0] _GEN_27912 = 6'h8 == state ? $signed(_GEN_307) : $signed(_GEN_27233); // @[digest.scala 81:19]
  wire [31:0] _GEN_27913 = 6'h8 == state ? $signed(_GEN_308) : $signed(_GEN_27234); // @[digest.scala 81:19]
  wire [31:0] _GEN_27914 = 6'h8 == state ? $signed(_GEN_309) : $signed(_GEN_27235); // @[digest.scala 81:19]
  wire [31:0] _GEN_27915 = 6'h8 == state ? $signed(_GEN_310) : $signed(_GEN_27236); // @[digest.scala 81:19]
  wire [31:0] _GEN_27916 = 6'h8 == state ? $signed(_GEN_311) : $signed(_GEN_27237); // @[digest.scala 81:19]
  wire [31:0] _GEN_27917 = 6'h8 == state ? $signed(_GEN_312) : $signed(_GEN_27238); // @[digest.scala 81:19]
  wire [31:0] _GEN_27918 = 6'h8 == state ? $signed(_GEN_313) : $signed(_GEN_27239); // @[digest.scala 81:19]
  wire [31:0] _GEN_27919 = 6'h8 == state ? $signed(_GEN_314) : $signed(_GEN_27240); // @[digest.scala 81:19]
  wire [31:0] _GEN_27920 = 6'h8 == state ? $signed(_GEN_315) : $signed(_GEN_27241); // @[digest.scala 81:19]
  wire [31:0] _GEN_27921 = 6'h8 == state ? $signed(_GEN_316) : $signed(_GEN_27242); // @[digest.scala 81:19]
  wire [31:0] _GEN_27922 = 6'h8 == state ? $signed(_GEN_317) : $signed(_GEN_27243); // @[digest.scala 81:19]
  wire [31:0] _GEN_27923 = 6'h8 == state ? $signed(_GEN_318) : $signed(_GEN_27244); // @[digest.scala 81:19]
  wire [31:0] _GEN_27924 = 6'h8 == state ? $signed(_GEN_319) : $signed(_GEN_27245); // @[digest.scala 81:19]
  wire [31:0] _GEN_27925 = 6'h8 == state ? $signed(_GEN_320) : $signed(_GEN_27246); // @[digest.scala 81:19]
  wire [5:0] _GEN_27926 = 6'h8 == state ? 6'h9 : _GEN_27247; // @[digest.scala 118:19 81:19]
  wire [31:0] _GEN_27927 = 6'h8 == state ? $signed(a) : $signed(_GEN_27248); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_27928 = 6'h8 == state ? $signed(b) : $signed(_GEN_27249); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_27929 = 6'h8 == state ? $signed(c) : $signed(_GEN_27250); // @[digest.scala 26:16 81:19]
  wire [31:0] _GEN_27930 = 6'h8 == state ? $signed(d) : $signed(_GEN_27251); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_27931 = 6'h8 == state ? $signed(e) : $signed(_GEN_27252); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_27932 = 6'h8 == state ? $signed(i) : $signed(_GEN_27253); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_27933 = 6'h8 == state ? $signed(olda) : $signed(_GEN_27254); // @[digest.scala 29:19 81:19]
  wire [31:0] _GEN_27934 = 6'h8 == state ? $signed(oldb) : $signed(_GEN_27255); // @[digest.scala 30:19 81:19]
  wire [31:0] _GEN_27935 = 6'h8 == state ? $signed(oldc) : $signed(_GEN_27256); // @[digest.scala 31:19 81:19]
  wire [31:0] _GEN_27936 = 6'h8 == state ? $signed(oldd) : $signed(_GEN_27257); // @[digest.scala 32:19 81:19]
  wire [31:0] _GEN_27937 = 6'h8 == state ? $signed(olde) : $signed(_GEN_27258); // @[digest.scala 33:19 81:19]
  wire [31:0] _GEN_27938 = 6'h8 == state ? $signed(j) : $signed(_GEN_27259); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_27939 = 6'h8 == state ? $signed(w_0) : $signed(_GEN_27260); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27940 = 6'h8 == state ? $signed(w_1) : $signed(_GEN_27261); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27941 = 6'h8 == state ? $signed(w_2) : $signed(_GEN_27262); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27942 = 6'h8 == state ? $signed(w_3) : $signed(_GEN_27263); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27943 = 6'h8 == state ? $signed(w_4) : $signed(_GEN_27264); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27944 = 6'h8 == state ? $signed(w_5) : $signed(_GEN_27265); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27945 = 6'h8 == state ? $signed(w_6) : $signed(_GEN_27266); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27946 = 6'h8 == state ? $signed(w_7) : $signed(_GEN_27267); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27947 = 6'h8 == state ? $signed(w_8) : $signed(_GEN_27268); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27948 = 6'h8 == state ? $signed(w_9) : $signed(_GEN_27269); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27949 = 6'h8 == state ? $signed(w_10) : $signed(_GEN_27270); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27950 = 6'h8 == state ? $signed(w_11) : $signed(_GEN_27271); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27951 = 6'h8 == state ? $signed(w_12) : $signed(_GEN_27272); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27952 = 6'h8 == state ? $signed(w_13) : $signed(_GEN_27273); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27953 = 6'h8 == state ? $signed(w_14) : $signed(_GEN_27274); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27954 = 6'h8 == state ? $signed(w_15) : $signed(_GEN_27275); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27955 = 6'h8 == state ? $signed(w_16) : $signed(_GEN_27276); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27956 = 6'h8 == state ? $signed(w_17) : $signed(_GEN_27277); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27957 = 6'h8 == state ? $signed(w_18) : $signed(_GEN_27278); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27958 = 6'h8 == state ? $signed(w_19) : $signed(_GEN_27279); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27959 = 6'h8 == state ? $signed(w_20) : $signed(_GEN_27280); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27960 = 6'h8 == state ? $signed(w_21) : $signed(_GEN_27281); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27961 = 6'h8 == state ? $signed(w_22) : $signed(_GEN_27282); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27962 = 6'h8 == state ? $signed(w_23) : $signed(_GEN_27283); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27963 = 6'h8 == state ? $signed(w_24) : $signed(_GEN_27284); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27964 = 6'h8 == state ? $signed(w_25) : $signed(_GEN_27285); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27965 = 6'h8 == state ? $signed(w_26) : $signed(_GEN_27286); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27966 = 6'h8 == state ? $signed(w_27) : $signed(_GEN_27287); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27967 = 6'h8 == state ? $signed(w_28) : $signed(_GEN_27288); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27968 = 6'h8 == state ? $signed(w_29) : $signed(_GEN_27289); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27969 = 6'h8 == state ? $signed(w_30) : $signed(_GEN_27290); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27970 = 6'h8 == state ? $signed(w_31) : $signed(_GEN_27291); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27971 = 6'h8 == state ? $signed(w_32) : $signed(_GEN_27292); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27972 = 6'h8 == state ? $signed(w_33) : $signed(_GEN_27293); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27973 = 6'h8 == state ? $signed(w_34) : $signed(_GEN_27294); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27974 = 6'h8 == state ? $signed(w_35) : $signed(_GEN_27295); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27975 = 6'h8 == state ? $signed(w_36) : $signed(_GEN_27296); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27976 = 6'h8 == state ? $signed(w_37) : $signed(_GEN_27297); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27977 = 6'h8 == state ? $signed(w_38) : $signed(_GEN_27298); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27978 = 6'h8 == state ? $signed(w_39) : $signed(_GEN_27299); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27979 = 6'h8 == state ? $signed(w_40) : $signed(_GEN_27300); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27980 = 6'h8 == state ? $signed(w_41) : $signed(_GEN_27301); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27981 = 6'h8 == state ? $signed(w_42) : $signed(_GEN_27302); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27982 = 6'h8 == state ? $signed(w_43) : $signed(_GEN_27303); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27983 = 6'h8 == state ? $signed(w_44) : $signed(_GEN_27304); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27984 = 6'h8 == state ? $signed(w_45) : $signed(_GEN_27305); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27985 = 6'h8 == state ? $signed(w_46) : $signed(_GEN_27306); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27986 = 6'h8 == state ? $signed(w_47) : $signed(_GEN_27307); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27987 = 6'h8 == state ? $signed(w_48) : $signed(_GEN_27308); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27988 = 6'h8 == state ? $signed(w_49) : $signed(_GEN_27309); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27989 = 6'h8 == state ? $signed(w_50) : $signed(_GEN_27310); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27990 = 6'h8 == state ? $signed(w_51) : $signed(_GEN_27311); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27991 = 6'h8 == state ? $signed(w_52) : $signed(_GEN_27312); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27992 = 6'h8 == state ? $signed(w_53) : $signed(_GEN_27313); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27993 = 6'h8 == state ? $signed(w_54) : $signed(_GEN_27314); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27994 = 6'h8 == state ? $signed(w_55) : $signed(_GEN_27315); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27995 = 6'h8 == state ? $signed(w_56) : $signed(_GEN_27316); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27996 = 6'h8 == state ? $signed(w_57) : $signed(_GEN_27317); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27997 = 6'h8 == state ? $signed(w_58) : $signed(_GEN_27318); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27998 = 6'h8 == state ? $signed(w_59) : $signed(_GEN_27319); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_27999 = 6'h8 == state ? $signed(w_60) : $signed(_GEN_27320); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28000 = 6'h8 == state ? $signed(w_61) : $signed(_GEN_27321); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28001 = 6'h8 == state ? $signed(w_62) : $signed(_GEN_27322); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28002 = 6'h8 == state ? $signed(w_63) : $signed(_GEN_27323); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28003 = 6'h8 == state ? $signed(w_64) : $signed(_GEN_27324); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28004 = 6'h8 == state ? $signed(w_65) : $signed(_GEN_27325); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28005 = 6'h8 == state ? $signed(w_66) : $signed(_GEN_27326); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28006 = 6'h8 == state ? $signed(w_67) : $signed(_GEN_27327); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28007 = 6'h8 == state ? $signed(w_68) : $signed(_GEN_27328); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28008 = 6'h8 == state ? $signed(w_69) : $signed(_GEN_27329); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28009 = 6'h8 == state ? $signed(w_70) : $signed(_GEN_27330); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28010 = 6'h8 == state ? $signed(w_71) : $signed(_GEN_27331); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28011 = 6'h8 == state ? $signed(w_72) : $signed(_GEN_27332); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28012 = 6'h8 == state ? $signed(w_73) : $signed(_GEN_27333); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28013 = 6'h8 == state ? $signed(w_74) : $signed(_GEN_27334); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28014 = 6'h8 == state ? $signed(w_75) : $signed(_GEN_27335); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28015 = 6'h8 == state ? $signed(w_76) : $signed(_GEN_27336); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28016 = 6'h8 == state ? $signed(w_77) : $signed(_GEN_27337); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28017 = 6'h8 == state ? $signed(w_78) : $signed(_GEN_27338); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28018 = 6'h8 == state ? $signed(w_79) : $signed(_GEN_27339); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28019 = 6'h8 == state ? $signed(temp) : $signed(_GEN_27340); // @[digest.scala 38:19 81:19]
  wire  _GEN_28020 = 6'h8 == state ? 1'h0 : _GEN_27341; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_28023 = 6'h8 == state ? $signed(t) : $signed(_GEN_27344); // @[digest.scala 35:16 81:19]
  wire  _GEN_28024 = 6'h8 == state ? 1'h0 : _GEN_27345; // @[digest.scala 81:19 48:24]
  wire  _GEN_28027 = 6'h8 == state ? 1'h0 : _GEN_27348; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_28111 = 6'h8 == state ? $signed(digest_0) : $signed(_GEN_27432); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28112 = 6'h8 == state ? $signed(digest_1) : $signed(_GEN_27433); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28113 = 6'h8 == state ? $signed(digest_2) : $signed(_GEN_27434); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28114 = 6'h8 == state ? $signed(digest_3) : $signed(_GEN_27435); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28115 = 6'h8 == state ? $signed(digest_4) : $signed(_GEN_27436); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28116 = 6'h8 == state ? $signed(digest_5) : $signed(_GEN_27437); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28117 = 6'h8 == state ? $signed(digest_6) : $signed(_GEN_27438); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28118 = 6'h8 == state ? $signed(digest_7) : $signed(_GEN_27439); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28119 = 6'h8 == state ? $signed(digest_8) : $signed(_GEN_27440); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28120 = 6'h8 == state ? $signed(digest_9) : $signed(_GEN_27441); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28121 = 6'h8 == state ? $signed(digest_10) : $signed(_GEN_27442); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28122 = 6'h8 == state ? $signed(digest_11) : $signed(_GEN_27443); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28123 = 6'h8 == state ? $signed(digest_12) : $signed(_GEN_27444); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28124 = 6'h8 == state ? $signed(digest_13) : $signed(_GEN_27445); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28125 = 6'h8 == state ? $signed(digest_14) : $signed(_GEN_27446); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28126 = 6'h8 == state ? $signed(digest_15) : $signed(_GEN_27447); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28127 = 6'h8 == state ? $signed(digest_16) : $signed(_GEN_27448); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28128 = 6'h8 == state ? $signed(digest_17) : $signed(_GEN_27449); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28129 = 6'h8 == state ? $signed(digest_18) : $signed(_GEN_27450); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28130 = 6'h8 == state ? $signed(digest_19) : $signed(_GEN_27451); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28131 = 6'h8 == state ? $signed(digest_20) : $signed(_GEN_27452); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28132 = 6'h8 == state ? $signed(digest_21) : $signed(_GEN_27453); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28133 = 6'h8 == state ? $signed(digest_22) : $signed(_GEN_27454); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28134 = 6'h8 == state ? $signed(digest_23) : $signed(_GEN_27455); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28135 = 6'h8 == state ? $signed(digest_24) : $signed(_GEN_27456); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28136 = 6'h8 == state ? $signed(digest_25) : $signed(_GEN_27457); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28137 = 6'h8 == state ? $signed(digest_26) : $signed(_GEN_27458); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28138 = 6'h8 == state ? $signed(digest_27) : $signed(_GEN_27459); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28139 = 6'h8 == state ? $signed(digest_28) : $signed(_GEN_27460); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28140 = 6'h8 == state ? $signed(digest_29) : $signed(_GEN_27461); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28141 = 6'h8 == state ? $signed(digest_30) : $signed(_GEN_27462); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28142 = 6'h8 == state ? $signed(digest_31) : $signed(_GEN_27463); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28143 = 6'h8 == state ? $signed(digest_32) : $signed(_GEN_27464); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28144 = 6'h8 == state ? $signed(digest_33) : $signed(_GEN_27465); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28145 = 6'h8 == state ? $signed(digest_34) : $signed(_GEN_27466); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28146 = 6'h8 == state ? $signed(digest_35) : $signed(_GEN_27467); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28147 = 6'h8 == state ? $signed(digest_36) : $signed(_GEN_27468); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28148 = 6'h8 == state ? $signed(digest_37) : $signed(_GEN_27469); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28149 = 6'h8 == state ? $signed(digest_38) : $signed(_GEN_27470); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28150 = 6'h8 == state ? $signed(digest_39) : $signed(_GEN_27471); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28151 = 6'h8 == state ? $signed(digest_40) : $signed(_GEN_27472); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28152 = 6'h8 == state ? $signed(digest_41) : $signed(_GEN_27473); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28153 = 6'h8 == state ? $signed(digest_42) : $signed(_GEN_27474); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28154 = 6'h8 == state ? $signed(digest_43) : $signed(_GEN_27475); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28155 = 6'h8 == state ? $signed(digest_44) : $signed(_GEN_27476); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28156 = 6'h8 == state ? $signed(digest_45) : $signed(_GEN_27477); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28157 = 6'h8 == state ? $signed(digest_46) : $signed(_GEN_27478); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28158 = 6'h8 == state ? $signed(digest_47) : $signed(_GEN_27479); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28159 = 6'h8 == state ? $signed(digest_48) : $signed(_GEN_27480); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28160 = 6'h8 == state ? $signed(digest_49) : $signed(_GEN_27481); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28161 = 6'h8 == state ? $signed(digest_50) : $signed(_GEN_27482); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28162 = 6'h8 == state ? $signed(digest_51) : $signed(_GEN_27483); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28163 = 6'h8 == state ? $signed(digest_52) : $signed(_GEN_27484); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28164 = 6'h8 == state ? $signed(digest_53) : $signed(_GEN_27485); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28165 = 6'h8 == state ? $signed(digest_54) : $signed(_GEN_27486); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28166 = 6'h8 == state ? $signed(digest_55) : $signed(_GEN_27487); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28167 = 6'h8 == state ? $signed(digest_56) : $signed(_GEN_27488); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28168 = 6'h8 == state ? $signed(digest_57) : $signed(_GEN_27489); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28169 = 6'h8 == state ? $signed(digest_58) : $signed(_GEN_27490); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28170 = 6'h8 == state ? $signed(digest_59) : $signed(_GEN_27491); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28171 = 6'h8 == state ? $signed(digest_60) : $signed(_GEN_27492); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28172 = 6'h8 == state ? $signed(digest_61) : $signed(_GEN_27493); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28173 = 6'h8 == state ? $signed(digest_62) : $signed(_GEN_27494); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28174 = 6'h8 == state ? $signed(digest_63) : $signed(_GEN_27495); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28175 = 6'h8 == state ? $signed(digest_64) : $signed(_GEN_27496); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28176 = 6'h8 == state ? $signed(digest_65) : $signed(_GEN_27497); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28177 = 6'h8 == state ? $signed(digest_66) : $signed(_GEN_27498); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28178 = 6'h8 == state ? $signed(digest_67) : $signed(_GEN_27499); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28179 = 6'h8 == state ? $signed(digest_68) : $signed(_GEN_27500); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28180 = 6'h8 == state ? $signed(digest_69) : $signed(_GEN_27501); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28181 = 6'h8 == state ? $signed(digest_70) : $signed(_GEN_27502); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28182 = 6'h8 == state ? $signed(digest_71) : $signed(_GEN_27503); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28183 = 6'h8 == state ? $signed(digest_72) : $signed(_GEN_27504); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28184 = 6'h8 == state ? $signed(digest_73) : $signed(_GEN_27505); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28185 = 6'h8 == state ? $signed(digest_74) : $signed(_GEN_27506); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28186 = 6'h8 == state ? $signed(digest_75) : $signed(_GEN_27507); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28187 = 6'h8 == state ? $signed(digest_76) : $signed(_GEN_27508); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28188 = 6'h8 == state ? $signed(digest_77) : $signed(_GEN_27509); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28189 = 6'h8 == state ? $signed(digest_78) : $signed(_GEN_27510); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28190 = 6'h8 == state ? $signed(digest_79) : $signed(_GEN_27511); // @[digest.scala 81:19 53:21]
  wire  _GEN_28192 = 6'h8 == state ? 1'h0 : _GEN_27513; // @[digest.scala 81:19 58:25]
  wire  _GEN_28275 = 6'h8 == state ? 1'h0 : _GEN_27596; // @[digest.scala 81:19 63:25]
  wire  _GEN_28358 = 6'h8 == state ? 1'h0 : _GEN_27679; // @[digest.scala 81:19 68:25]
  wire  _GEN_28441 = 6'h8 == state ? 1'h0 : _GEN_27762; // @[digest.scala 81:19 73:25]
  wire  _GEN_28524 = 6'h8 == state ? 1'h0 : _GEN_27845; // @[digest.scala 81:19 78:25]
  wire [62:0] _GEN_28525 = 6'h7 == state ? $signed(_temp_T_17) : $signed({{31{_GEN_28019[31]}},_GEN_28019}); // @[digest.scala 113:18 81:19]
  wire [5:0] _GEN_28526 = 6'h7 == state ? 6'h8 : _GEN_27926; // @[digest.scala 114:19 81:19]
  wire [31:0] _GEN_28527 = 6'h7 == state ? $signed(blks_0) : $signed(_GEN_27846); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28528 = 6'h7 == state ? $signed(blks_1) : $signed(_GEN_27847); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28529 = 6'h7 == state ? $signed(blks_2) : $signed(_GEN_27848); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28530 = 6'h7 == state ? $signed(blks_3) : $signed(_GEN_27849); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28531 = 6'h7 == state ? $signed(blks_4) : $signed(_GEN_27850); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28532 = 6'h7 == state ? $signed(blks_5) : $signed(_GEN_27851); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28533 = 6'h7 == state ? $signed(blks_6) : $signed(_GEN_27852); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28534 = 6'h7 == state ? $signed(blks_7) : $signed(_GEN_27853); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28535 = 6'h7 == state ? $signed(blks_8) : $signed(_GEN_27854); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28536 = 6'h7 == state ? $signed(blks_9) : $signed(_GEN_27855); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28537 = 6'h7 == state ? $signed(blks_10) : $signed(_GEN_27856); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28538 = 6'h7 == state ? $signed(blks_11) : $signed(_GEN_27857); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28539 = 6'h7 == state ? $signed(blks_12) : $signed(_GEN_27858); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28540 = 6'h7 == state ? $signed(blks_13) : $signed(_GEN_27859); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28541 = 6'h7 == state ? $signed(blks_14) : $signed(_GEN_27860); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28542 = 6'h7 == state ? $signed(blks_15) : $signed(_GEN_27861); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28543 = 6'h7 == state ? $signed(blks_16) : $signed(_GEN_27862); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28544 = 6'h7 == state ? $signed(blks_17) : $signed(_GEN_27863); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28545 = 6'h7 == state ? $signed(blks_18) : $signed(_GEN_27864); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28546 = 6'h7 == state ? $signed(blks_19) : $signed(_GEN_27865); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28547 = 6'h7 == state ? $signed(blks_20) : $signed(_GEN_27866); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28548 = 6'h7 == state ? $signed(blks_21) : $signed(_GEN_27867); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28549 = 6'h7 == state ? $signed(blks_22) : $signed(_GEN_27868); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28550 = 6'h7 == state ? $signed(blks_23) : $signed(_GEN_27869); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28551 = 6'h7 == state ? $signed(blks_24) : $signed(_GEN_27870); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28552 = 6'h7 == state ? $signed(blks_25) : $signed(_GEN_27871); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28553 = 6'h7 == state ? $signed(blks_26) : $signed(_GEN_27872); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28554 = 6'h7 == state ? $signed(blks_27) : $signed(_GEN_27873); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28555 = 6'h7 == state ? $signed(blks_28) : $signed(_GEN_27874); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28556 = 6'h7 == state ? $signed(blks_29) : $signed(_GEN_27875); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28557 = 6'h7 == state ? $signed(blks_30) : $signed(_GEN_27876); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28558 = 6'h7 == state ? $signed(blks_31) : $signed(_GEN_27877); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28559 = 6'h7 == state ? $signed(blks_32) : $signed(_GEN_27878); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28560 = 6'h7 == state ? $signed(blks_33) : $signed(_GEN_27879); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28561 = 6'h7 == state ? $signed(blks_34) : $signed(_GEN_27880); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28562 = 6'h7 == state ? $signed(blks_35) : $signed(_GEN_27881); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28563 = 6'h7 == state ? $signed(blks_36) : $signed(_GEN_27882); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28564 = 6'h7 == state ? $signed(blks_37) : $signed(_GEN_27883); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28565 = 6'h7 == state ? $signed(blks_38) : $signed(_GEN_27884); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28566 = 6'h7 == state ? $signed(blks_39) : $signed(_GEN_27885); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28567 = 6'h7 == state ? $signed(blks_40) : $signed(_GEN_27886); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28568 = 6'h7 == state ? $signed(blks_41) : $signed(_GEN_27887); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28569 = 6'h7 == state ? $signed(blks_42) : $signed(_GEN_27888); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28570 = 6'h7 == state ? $signed(blks_43) : $signed(_GEN_27889); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28571 = 6'h7 == state ? $signed(blks_44) : $signed(_GEN_27890); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28572 = 6'h7 == state ? $signed(blks_45) : $signed(_GEN_27891); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28573 = 6'h7 == state ? $signed(blks_46) : $signed(_GEN_27892); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28574 = 6'h7 == state ? $signed(blks_47) : $signed(_GEN_27893); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28575 = 6'h7 == state ? $signed(blks_48) : $signed(_GEN_27894); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28576 = 6'h7 == state ? $signed(blks_49) : $signed(_GEN_27895); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28577 = 6'h7 == state ? $signed(blks_50) : $signed(_GEN_27896); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28578 = 6'h7 == state ? $signed(blks_51) : $signed(_GEN_27897); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28579 = 6'h7 == state ? $signed(blks_52) : $signed(_GEN_27898); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28580 = 6'h7 == state ? $signed(blks_53) : $signed(_GEN_27899); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28581 = 6'h7 == state ? $signed(blks_54) : $signed(_GEN_27900); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28582 = 6'h7 == state ? $signed(blks_55) : $signed(_GEN_27901); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28583 = 6'h7 == state ? $signed(blks_56) : $signed(_GEN_27902); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28584 = 6'h7 == state ? $signed(blks_57) : $signed(_GEN_27903); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28585 = 6'h7 == state ? $signed(blks_58) : $signed(_GEN_27904); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28586 = 6'h7 == state ? $signed(blks_59) : $signed(_GEN_27905); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28587 = 6'h7 == state ? $signed(blks_60) : $signed(_GEN_27906); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28588 = 6'h7 == state ? $signed(blks_61) : $signed(_GEN_27907); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28589 = 6'h7 == state ? $signed(blks_62) : $signed(_GEN_27908); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28590 = 6'h7 == state ? $signed(blks_63) : $signed(_GEN_27909); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28591 = 6'h7 == state ? $signed(blks_64) : $signed(_GEN_27910); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28592 = 6'h7 == state ? $signed(blks_65) : $signed(_GEN_27911); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28593 = 6'h7 == state ? $signed(blks_66) : $signed(_GEN_27912); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28594 = 6'h7 == state ? $signed(blks_67) : $signed(_GEN_27913); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28595 = 6'h7 == state ? $signed(blks_68) : $signed(_GEN_27914); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28596 = 6'h7 == state ? $signed(blks_69) : $signed(_GEN_27915); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28597 = 6'h7 == state ? $signed(blks_70) : $signed(_GEN_27916); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28598 = 6'h7 == state ? $signed(blks_71) : $signed(_GEN_27917); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28599 = 6'h7 == state ? $signed(blks_72) : $signed(_GEN_27918); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28600 = 6'h7 == state ? $signed(blks_73) : $signed(_GEN_27919); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28601 = 6'h7 == state ? $signed(blks_74) : $signed(_GEN_27920); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28602 = 6'h7 == state ? $signed(blks_75) : $signed(_GEN_27921); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28603 = 6'h7 == state ? $signed(blks_76) : $signed(_GEN_27922); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28604 = 6'h7 == state ? $signed(blks_77) : $signed(_GEN_27923); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28605 = 6'h7 == state ? $signed(blks_78) : $signed(_GEN_27924); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28606 = 6'h7 == state ? $signed(blks_79) : $signed(_GEN_27925); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_28607 = 6'h7 == state ? $signed(a) : $signed(_GEN_27927); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_28608 = 6'h7 == state ? $signed(b) : $signed(_GEN_27928); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_28609 = 6'h7 == state ? $signed(c) : $signed(_GEN_27929); // @[digest.scala 26:16 81:19]
  wire [31:0] _GEN_28610 = 6'h7 == state ? $signed(d) : $signed(_GEN_27930); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_28611 = 6'h7 == state ? $signed(e) : $signed(_GEN_27931); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_28612 = 6'h7 == state ? $signed(i) : $signed(_GEN_27932); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_28613 = 6'h7 == state ? $signed(olda) : $signed(_GEN_27933); // @[digest.scala 29:19 81:19]
  wire [31:0] _GEN_28614 = 6'h7 == state ? $signed(oldb) : $signed(_GEN_27934); // @[digest.scala 30:19 81:19]
  wire [31:0] _GEN_28615 = 6'h7 == state ? $signed(oldc) : $signed(_GEN_27935); // @[digest.scala 31:19 81:19]
  wire [31:0] _GEN_28616 = 6'h7 == state ? $signed(oldd) : $signed(_GEN_27936); // @[digest.scala 32:19 81:19]
  wire [31:0] _GEN_28617 = 6'h7 == state ? $signed(olde) : $signed(_GEN_27937); // @[digest.scala 33:19 81:19]
  wire [31:0] _GEN_28618 = 6'h7 == state ? $signed(j) : $signed(_GEN_27938); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_28619 = 6'h7 == state ? $signed(w_0) : $signed(_GEN_27939); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28620 = 6'h7 == state ? $signed(w_1) : $signed(_GEN_27940); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28621 = 6'h7 == state ? $signed(w_2) : $signed(_GEN_27941); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28622 = 6'h7 == state ? $signed(w_3) : $signed(_GEN_27942); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28623 = 6'h7 == state ? $signed(w_4) : $signed(_GEN_27943); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28624 = 6'h7 == state ? $signed(w_5) : $signed(_GEN_27944); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28625 = 6'h7 == state ? $signed(w_6) : $signed(_GEN_27945); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28626 = 6'h7 == state ? $signed(w_7) : $signed(_GEN_27946); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28627 = 6'h7 == state ? $signed(w_8) : $signed(_GEN_27947); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28628 = 6'h7 == state ? $signed(w_9) : $signed(_GEN_27948); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28629 = 6'h7 == state ? $signed(w_10) : $signed(_GEN_27949); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28630 = 6'h7 == state ? $signed(w_11) : $signed(_GEN_27950); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28631 = 6'h7 == state ? $signed(w_12) : $signed(_GEN_27951); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28632 = 6'h7 == state ? $signed(w_13) : $signed(_GEN_27952); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28633 = 6'h7 == state ? $signed(w_14) : $signed(_GEN_27953); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28634 = 6'h7 == state ? $signed(w_15) : $signed(_GEN_27954); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28635 = 6'h7 == state ? $signed(w_16) : $signed(_GEN_27955); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28636 = 6'h7 == state ? $signed(w_17) : $signed(_GEN_27956); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28637 = 6'h7 == state ? $signed(w_18) : $signed(_GEN_27957); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28638 = 6'h7 == state ? $signed(w_19) : $signed(_GEN_27958); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28639 = 6'h7 == state ? $signed(w_20) : $signed(_GEN_27959); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28640 = 6'h7 == state ? $signed(w_21) : $signed(_GEN_27960); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28641 = 6'h7 == state ? $signed(w_22) : $signed(_GEN_27961); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28642 = 6'h7 == state ? $signed(w_23) : $signed(_GEN_27962); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28643 = 6'h7 == state ? $signed(w_24) : $signed(_GEN_27963); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28644 = 6'h7 == state ? $signed(w_25) : $signed(_GEN_27964); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28645 = 6'h7 == state ? $signed(w_26) : $signed(_GEN_27965); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28646 = 6'h7 == state ? $signed(w_27) : $signed(_GEN_27966); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28647 = 6'h7 == state ? $signed(w_28) : $signed(_GEN_27967); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28648 = 6'h7 == state ? $signed(w_29) : $signed(_GEN_27968); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28649 = 6'h7 == state ? $signed(w_30) : $signed(_GEN_27969); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28650 = 6'h7 == state ? $signed(w_31) : $signed(_GEN_27970); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28651 = 6'h7 == state ? $signed(w_32) : $signed(_GEN_27971); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28652 = 6'h7 == state ? $signed(w_33) : $signed(_GEN_27972); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28653 = 6'h7 == state ? $signed(w_34) : $signed(_GEN_27973); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28654 = 6'h7 == state ? $signed(w_35) : $signed(_GEN_27974); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28655 = 6'h7 == state ? $signed(w_36) : $signed(_GEN_27975); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28656 = 6'h7 == state ? $signed(w_37) : $signed(_GEN_27976); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28657 = 6'h7 == state ? $signed(w_38) : $signed(_GEN_27977); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28658 = 6'h7 == state ? $signed(w_39) : $signed(_GEN_27978); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28659 = 6'h7 == state ? $signed(w_40) : $signed(_GEN_27979); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28660 = 6'h7 == state ? $signed(w_41) : $signed(_GEN_27980); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28661 = 6'h7 == state ? $signed(w_42) : $signed(_GEN_27981); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28662 = 6'h7 == state ? $signed(w_43) : $signed(_GEN_27982); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28663 = 6'h7 == state ? $signed(w_44) : $signed(_GEN_27983); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28664 = 6'h7 == state ? $signed(w_45) : $signed(_GEN_27984); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28665 = 6'h7 == state ? $signed(w_46) : $signed(_GEN_27985); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28666 = 6'h7 == state ? $signed(w_47) : $signed(_GEN_27986); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28667 = 6'h7 == state ? $signed(w_48) : $signed(_GEN_27987); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28668 = 6'h7 == state ? $signed(w_49) : $signed(_GEN_27988); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28669 = 6'h7 == state ? $signed(w_50) : $signed(_GEN_27989); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28670 = 6'h7 == state ? $signed(w_51) : $signed(_GEN_27990); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28671 = 6'h7 == state ? $signed(w_52) : $signed(_GEN_27991); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28672 = 6'h7 == state ? $signed(w_53) : $signed(_GEN_27992); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28673 = 6'h7 == state ? $signed(w_54) : $signed(_GEN_27993); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28674 = 6'h7 == state ? $signed(w_55) : $signed(_GEN_27994); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28675 = 6'h7 == state ? $signed(w_56) : $signed(_GEN_27995); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28676 = 6'h7 == state ? $signed(w_57) : $signed(_GEN_27996); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28677 = 6'h7 == state ? $signed(w_58) : $signed(_GEN_27997); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28678 = 6'h7 == state ? $signed(w_59) : $signed(_GEN_27998); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28679 = 6'h7 == state ? $signed(w_60) : $signed(_GEN_27999); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28680 = 6'h7 == state ? $signed(w_61) : $signed(_GEN_28000); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28681 = 6'h7 == state ? $signed(w_62) : $signed(_GEN_28001); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28682 = 6'h7 == state ? $signed(w_63) : $signed(_GEN_28002); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28683 = 6'h7 == state ? $signed(w_64) : $signed(_GEN_28003); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28684 = 6'h7 == state ? $signed(w_65) : $signed(_GEN_28004); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28685 = 6'h7 == state ? $signed(w_66) : $signed(_GEN_28005); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28686 = 6'h7 == state ? $signed(w_67) : $signed(_GEN_28006); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28687 = 6'h7 == state ? $signed(w_68) : $signed(_GEN_28007); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28688 = 6'h7 == state ? $signed(w_69) : $signed(_GEN_28008); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28689 = 6'h7 == state ? $signed(w_70) : $signed(_GEN_28009); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28690 = 6'h7 == state ? $signed(w_71) : $signed(_GEN_28010); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28691 = 6'h7 == state ? $signed(w_72) : $signed(_GEN_28011); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28692 = 6'h7 == state ? $signed(w_73) : $signed(_GEN_28012); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28693 = 6'h7 == state ? $signed(w_74) : $signed(_GEN_28013); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28694 = 6'h7 == state ? $signed(w_75) : $signed(_GEN_28014); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28695 = 6'h7 == state ? $signed(w_76) : $signed(_GEN_28015); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28696 = 6'h7 == state ? $signed(w_77) : $signed(_GEN_28016); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28697 = 6'h7 == state ? $signed(w_78) : $signed(_GEN_28017); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_28698 = 6'h7 == state ? $signed(w_79) : $signed(_GEN_28018); // @[digest.scala 40:16 81:19]
  wire  _GEN_28699 = 6'h7 == state ? 1'h0 : _GEN_28020; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_28702 = 6'h7 == state ? $signed(t) : $signed(_GEN_28023); // @[digest.scala 35:16 81:19]
  wire  _GEN_28703 = 6'h7 == state ? 1'h0 : _GEN_28024; // @[digest.scala 81:19 48:24]
  wire  _GEN_28706 = 6'h7 == state ? 1'h0 : _GEN_28027; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_28790 = 6'h7 == state ? $signed(digest_0) : $signed(_GEN_28111); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28791 = 6'h7 == state ? $signed(digest_1) : $signed(_GEN_28112); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28792 = 6'h7 == state ? $signed(digest_2) : $signed(_GEN_28113); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28793 = 6'h7 == state ? $signed(digest_3) : $signed(_GEN_28114); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28794 = 6'h7 == state ? $signed(digest_4) : $signed(_GEN_28115); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28795 = 6'h7 == state ? $signed(digest_5) : $signed(_GEN_28116); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28796 = 6'h7 == state ? $signed(digest_6) : $signed(_GEN_28117); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28797 = 6'h7 == state ? $signed(digest_7) : $signed(_GEN_28118); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28798 = 6'h7 == state ? $signed(digest_8) : $signed(_GEN_28119); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28799 = 6'h7 == state ? $signed(digest_9) : $signed(_GEN_28120); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28800 = 6'h7 == state ? $signed(digest_10) : $signed(_GEN_28121); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28801 = 6'h7 == state ? $signed(digest_11) : $signed(_GEN_28122); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28802 = 6'h7 == state ? $signed(digest_12) : $signed(_GEN_28123); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28803 = 6'h7 == state ? $signed(digest_13) : $signed(_GEN_28124); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28804 = 6'h7 == state ? $signed(digest_14) : $signed(_GEN_28125); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28805 = 6'h7 == state ? $signed(digest_15) : $signed(_GEN_28126); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28806 = 6'h7 == state ? $signed(digest_16) : $signed(_GEN_28127); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28807 = 6'h7 == state ? $signed(digest_17) : $signed(_GEN_28128); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28808 = 6'h7 == state ? $signed(digest_18) : $signed(_GEN_28129); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28809 = 6'h7 == state ? $signed(digest_19) : $signed(_GEN_28130); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28810 = 6'h7 == state ? $signed(digest_20) : $signed(_GEN_28131); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28811 = 6'h7 == state ? $signed(digest_21) : $signed(_GEN_28132); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28812 = 6'h7 == state ? $signed(digest_22) : $signed(_GEN_28133); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28813 = 6'h7 == state ? $signed(digest_23) : $signed(_GEN_28134); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28814 = 6'h7 == state ? $signed(digest_24) : $signed(_GEN_28135); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28815 = 6'h7 == state ? $signed(digest_25) : $signed(_GEN_28136); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28816 = 6'h7 == state ? $signed(digest_26) : $signed(_GEN_28137); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28817 = 6'h7 == state ? $signed(digest_27) : $signed(_GEN_28138); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28818 = 6'h7 == state ? $signed(digest_28) : $signed(_GEN_28139); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28819 = 6'h7 == state ? $signed(digest_29) : $signed(_GEN_28140); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28820 = 6'h7 == state ? $signed(digest_30) : $signed(_GEN_28141); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28821 = 6'h7 == state ? $signed(digest_31) : $signed(_GEN_28142); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28822 = 6'h7 == state ? $signed(digest_32) : $signed(_GEN_28143); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28823 = 6'h7 == state ? $signed(digest_33) : $signed(_GEN_28144); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28824 = 6'h7 == state ? $signed(digest_34) : $signed(_GEN_28145); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28825 = 6'h7 == state ? $signed(digest_35) : $signed(_GEN_28146); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28826 = 6'h7 == state ? $signed(digest_36) : $signed(_GEN_28147); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28827 = 6'h7 == state ? $signed(digest_37) : $signed(_GEN_28148); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28828 = 6'h7 == state ? $signed(digest_38) : $signed(_GEN_28149); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28829 = 6'h7 == state ? $signed(digest_39) : $signed(_GEN_28150); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28830 = 6'h7 == state ? $signed(digest_40) : $signed(_GEN_28151); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28831 = 6'h7 == state ? $signed(digest_41) : $signed(_GEN_28152); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28832 = 6'h7 == state ? $signed(digest_42) : $signed(_GEN_28153); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28833 = 6'h7 == state ? $signed(digest_43) : $signed(_GEN_28154); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28834 = 6'h7 == state ? $signed(digest_44) : $signed(_GEN_28155); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28835 = 6'h7 == state ? $signed(digest_45) : $signed(_GEN_28156); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28836 = 6'h7 == state ? $signed(digest_46) : $signed(_GEN_28157); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28837 = 6'h7 == state ? $signed(digest_47) : $signed(_GEN_28158); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28838 = 6'h7 == state ? $signed(digest_48) : $signed(_GEN_28159); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28839 = 6'h7 == state ? $signed(digest_49) : $signed(_GEN_28160); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28840 = 6'h7 == state ? $signed(digest_50) : $signed(_GEN_28161); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28841 = 6'h7 == state ? $signed(digest_51) : $signed(_GEN_28162); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28842 = 6'h7 == state ? $signed(digest_52) : $signed(_GEN_28163); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28843 = 6'h7 == state ? $signed(digest_53) : $signed(_GEN_28164); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28844 = 6'h7 == state ? $signed(digest_54) : $signed(_GEN_28165); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28845 = 6'h7 == state ? $signed(digest_55) : $signed(_GEN_28166); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28846 = 6'h7 == state ? $signed(digest_56) : $signed(_GEN_28167); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28847 = 6'h7 == state ? $signed(digest_57) : $signed(_GEN_28168); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28848 = 6'h7 == state ? $signed(digest_58) : $signed(_GEN_28169); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28849 = 6'h7 == state ? $signed(digest_59) : $signed(_GEN_28170); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28850 = 6'h7 == state ? $signed(digest_60) : $signed(_GEN_28171); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28851 = 6'h7 == state ? $signed(digest_61) : $signed(_GEN_28172); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28852 = 6'h7 == state ? $signed(digest_62) : $signed(_GEN_28173); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28853 = 6'h7 == state ? $signed(digest_63) : $signed(_GEN_28174); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28854 = 6'h7 == state ? $signed(digest_64) : $signed(_GEN_28175); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28855 = 6'h7 == state ? $signed(digest_65) : $signed(_GEN_28176); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28856 = 6'h7 == state ? $signed(digest_66) : $signed(_GEN_28177); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28857 = 6'h7 == state ? $signed(digest_67) : $signed(_GEN_28178); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28858 = 6'h7 == state ? $signed(digest_68) : $signed(_GEN_28179); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28859 = 6'h7 == state ? $signed(digest_69) : $signed(_GEN_28180); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28860 = 6'h7 == state ? $signed(digest_70) : $signed(_GEN_28181); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28861 = 6'h7 == state ? $signed(digest_71) : $signed(_GEN_28182); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28862 = 6'h7 == state ? $signed(digest_72) : $signed(_GEN_28183); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28863 = 6'h7 == state ? $signed(digest_73) : $signed(_GEN_28184); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28864 = 6'h7 == state ? $signed(digest_74) : $signed(_GEN_28185); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28865 = 6'h7 == state ? $signed(digest_75) : $signed(_GEN_28186); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28866 = 6'h7 == state ? $signed(digest_76) : $signed(_GEN_28187); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28867 = 6'h7 == state ? $signed(digest_77) : $signed(_GEN_28188); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28868 = 6'h7 == state ? $signed(digest_78) : $signed(_GEN_28189); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_28869 = 6'h7 == state ? $signed(digest_79) : $signed(_GEN_28190); // @[digest.scala 81:19 53:21]
  wire  _GEN_28871 = 6'h7 == state ? 1'h0 : _GEN_28192; // @[digest.scala 81:19 58:25]
  wire  _GEN_28954 = 6'h7 == state ? 1'h0 : _GEN_28275; // @[digest.scala 81:19 63:25]
  wire  _GEN_29037 = 6'h7 == state ? 1'h0 : _GEN_28358; // @[digest.scala 81:19 68:25]
  wire  _GEN_29120 = 6'h7 == state ? 1'h0 : _GEN_28441; // @[digest.scala 81:19 73:25]
  wire  _GEN_29203 = 6'h7 == state ? 1'h0 : _GEN_28524; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_29204 = 6'h6 == state ? $signed(_i_T_2) : $signed(_GEN_28612); // @[digest.scala 109:15 81:19]
  wire [5:0] _GEN_29205 = 6'h6 == state ? 6'h3 : _GEN_28526; // @[digest.scala 110:19 81:19]
  wire [62:0] _GEN_29206 = 6'h6 == state ? $signed({{31{temp[31]}},temp}) : $signed(_GEN_28525); // @[digest.scala 38:19 81:19]
  wire [31:0] _GEN_29207 = 6'h6 == state ? $signed(blks_0) : $signed(_GEN_28527); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29208 = 6'h6 == state ? $signed(blks_1) : $signed(_GEN_28528); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29209 = 6'h6 == state ? $signed(blks_2) : $signed(_GEN_28529); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29210 = 6'h6 == state ? $signed(blks_3) : $signed(_GEN_28530); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29211 = 6'h6 == state ? $signed(blks_4) : $signed(_GEN_28531); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29212 = 6'h6 == state ? $signed(blks_5) : $signed(_GEN_28532); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29213 = 6'h6 == state ? $signed(blks_6) : $signed(_GEN_28533); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29214 = 6'h6 == state ? $signed(blks_7) : $signed(_GEN_28534); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29215 = 6'h6 == state ? $signed(blks_8) : $signed(_GEN_28535); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29216 = 6'h6 == state ? $signed(blks_9) : $signed(_GEN_28536); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29217 = 6'h6 == state ? $signed(blks_10) : $signed(_GEN_28537); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29218 = 6'h6 == state ? $signed(blks_11) : $signed(_GEN_28538); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29219 = 6'h6 == state ? $signed(blks_12) : $signed(_GEN_28539); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29220 = 6'h6 == state ? $signed(blks_13) : $signed(_GEN_28540); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29221 = 6'h6 == state ? $signed(blks_14) : $signed(_GEN_28541); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29222 = 6'h6 == state ? $signed(blks_15) : $signed(_GEN_28542); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29223 = 6'h6 == state ? $signed(blks_16) : $signed(_GEN_28543); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29224 = 6'h6 == state ? $signed(blks_17) : $signed(_GEN_28544); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29225 = 6'h6 == state ? $signed(blks_18) : $signed(_GEN_28545); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29226 = 6'h6 == state ? $signed(blks_19) : $signed(_GEN_28546); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29227 = 6'h6 == state ? $signed(blks_20) : $signed(_GEN_28547); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29228 = 6'h6 == state ? $signed(blks_21) : $signed(_GEN_28548); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29229 = 6'h6 == state ? $signed(blks_22) : $signed(_GEN_28549); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29230 = 6'h6 == state ? $signed(blks_23) : $signed(_GEN_28550); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29231 = 6'h6 == state ? $signed(blks_24) : $signed(_GEN_28551); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29232 = 6'h6 == state ? $signed(blks_25) : $signed(_GEN_28552); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29233 = 6'h6 == state ? $signed(blks_26) : $signed(_GEN_28553); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29234 = 6'h6 == state ? $signed(blks_27) : $signed(_GEN_28554); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29235 = 6'h6 == state ? $signed(blks_28) : $signed(_GEN_28555); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29236 = 6'h6 == state ? $signed(blks_29) : $signed(_GEN_28556); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29237 = 6'h6 == state ? $signed(blks_30) : $signed(_GEN_28557); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29238 = 6'h6 == state ? $signed(blks_31) : $signed(_GEN_28558); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29239 = 6'h6 == state ? $signed(blks_32) : $signed(_GEN_28559); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29240 = 6'h6 == state ? $signed(blks_33) : $signed(_GEN_28560); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29241 = 6'h6 == state ? $signed(blks_34) : $signed(_GEN_28561); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29242 = 6'h6 == state ? $signed(blks_35) : $signed(_GEN_28562); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29243 = 6'h6 == state ? $signed(blks_36) : $signed(_GEN_28563); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29244 = 6'h6 == state ? $signed(blks_37) : $signed(_GEN_28564); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29245 = 6'h6 == state ? $signed(blks_38) : $signed(_GEN_28565); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29246 = 6'h6 == state ? $signed(blks_39) : $signed(_GEN_28566); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29247 = 6'h6 == state ? $signed(blks_40) : $signed(_GEN_28567); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29248 = 6'h6 == state ? $signed(blks_41) : $signed(_GEN_28568); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29249 = 6'h6 == state ? $signed(blks_42) : $signed(_GEN_28569); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29250 = 6'h6 == state ? $signed(blks_43) : $signed(_GEN_28570); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29251 = 6'h6 == state ? $signed(blks_44) : $signed(_GEN_28571); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29252 = 6'h6 == state ? $signed(blks_45) : $signed(_GEN_28572); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29253 = 6'h6 == state ? $signed(blks_46) : $signed(_GEN_28573); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29254 = 6'h6 == state ? $signed(blks_47) : $signed(_GEN_28574); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29255 = 6'h6 == state ? $signed(blks_48) : $signed(_GEN_28575); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29256 = 6'h6 == state ? $signed(blks_49) : $signed(_GEN_28576); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29257 = 6'h6 == state ? $signed(blks_50) : $signed(_GEN_28577); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29258 = 6'h6 == state ? $signed(blks_51) : $signed(_GEN_28578); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29259 = 6'h6 == state ? $signed(blks_52) : $signed(_GEN_28579); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29260 = 6'h6 == state ? $signed(blks_53) : $signed(_GEN_28580); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29261 = 6'h6 == state ? $signed(blks_54) : $signed(_GEN_28581); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29262 = 6'h6 == state ? $signed(blks_55) : $signed(_GEN_28582); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29263 = 6'h6 == state ? $signed(blks_56) : $signed(_GEN_28583); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29264 = 6'h6 == state ? $signed(blks_57) : $signed(_GEN_28584); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29265 = 6'h6 == state ? $signed(blks_58) : $signed(_GEN_28585); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29266 = 6'h6 == state ? $signed(blks_59) : $signed(_GEN_28586); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29267 = 6'h6 == state ? $signed(blks_60) : $signed(_GEN_28587); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29268 = 6'h6 == state ? $signed(blks_61) : $signed(_GEN_28588); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29269 = 6'h6 == state ? $signed(blks_62) : $signed(_GEN_28589); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29270 = 6'h6 == state ? $signed(blks_63) : $signed(_GEN_28590); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29271 = 6'h6 == state ? $signed(blks_64) : $signed(_GEN_28591); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29272 = 6'h6 == state ? $signed(blks_65) : $signed(_GEN_28592); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29273 = 6'h6 == state ? $signed(blks_66) : $signed(_GEN_28593); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29274 = 6'h6 == state ? $signed(blks_67) : $signed(_GEN_28594); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29275 = 6'h6 == state ? $signed(blks_68) : $signed(_GEN_28595); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29276 = 6'h6 == state ? $signed(blks_69) : $signed(_GEN_28596); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29277 = 6'h6 == state ? $signed(blks_70) : $signed(_GEN_28597); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29278 = 6'h6 == state ? $signed(blks_71) : $signed(_GEN_28598); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29279 = 6'h6 == state ? $signed(blks_72) : $signed(_GEN_28599); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29280 = 6'h6 == state ? $signed(blks_73) : $signed(_GEN_28600); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29281 = 6'h6 == state ? $signed(blks_74) : $signed(_GEN_28601); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29282 = 6'h6 == state ? $signed(blks_75) : $signed(_GEN_28602); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29283 = 6'h6 == state ? $signed(blks_76) : $signed(_GEN_28603); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29284 = 6'h6 == state ? $signed(blks_77) : $signed(_GEN_28604); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29285 = 6'h6 == state ? $signed(blks_78) : $signed(_GEN_28605); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29286 = 6'h6 == state ? $signed(blks_79) : $signed(_GEN_28606); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_29287 = 6'h6 == state ? $signed(a) : $signed(_GEN_28607); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_29288 = 6'h6 == state ? $signed(b) : $signed(_GEN_28608); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_29289 = 6'h6 == state ? $signed(c) : $signed(_GEN_28609); // @[digest.scala 26:16 81:19]
  wire [31:0] _GEN_29290 = 6'h6 == state ? $signed(d) : $signed(_GEN_28610); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_29291 = 6'h6 == state ? $signed(e) : $signed(_GEN_28611); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_29292 = 6'h6 == state ? $signed(olda) : $signed(_GEN_28613); // @[digest.scala 29:19 81:19]
  wire [31:0] _GEN_29293 = 6'h6 == state ? $signed(oldb) : $signed(_GEN_28614); // @[digest.scala 30:19 81:19]
  wire [31:0] _GEN_29294 = 6'h6 == state ? $signed(oldc) : $signed(_GEN_28615); // @[digest.scala 31:19 81:19]
  wire [31:0] _GEN_29295 = 6'h6 == state ? $signed(oldd) : $signed(_GEN_28616); // @[digest.scala 32:19 81:19]
  wire [31:0] _GEN_29296 = 6'h6 == state ? $signed(olde) : $signed(_GEN_28617); // @[digest.scala 33:19 81:19]
  wire [31:0] _GEN_29297 = 6'h6 == state ? $signed(j) : $signed(_GEN_28618); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_29298 = 6'h6 == state ? $signed(w_0) : $signed(_GEN_28619); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29299 = 6'h6 == state ? $signed(w_1) : $signed(_GEN_28620); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29300 = 6'h6 == state ? $signed(w_2) : $signed(_GEN_28621); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29301 = 6'h6 == state ? $signed(w_3) : $signed(_GEN_28622); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29302 = 6'h6 == state ? $signed(w_4) : $signed(_GEN_28623); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29303 = 6'h6 == state ? $signed(w_5) : $signed(_GEN_28624); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29304 = 6'h6 == state ? $signed(w_6) : $signed(_GEN_28625); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29305 = 6'h6 == state ? $signed(w_7) : $signed(_GEN_28626); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29306 = 6'h6 == state ? $signed(w_8) : $signed(_GEN_28627); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29307 = 6'h6 == state ? $signed(w_9) : $signed(_GEN_28628); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29308 = 6'h6 == state ? $signed(w_10) : $signed(_GEN_28629); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29309 = 6'h6 == state ? $signed(w_11) : $signed(_GEN_28630); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29310 = 6'h6 == state ? $signed(w_12) : $signed(_GEN_28631); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29311 = 6'h6 == state ? $signed(w_13) : $signed(_GEN_28632); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29312 = 6'h6 == state ? $signed(w_14) : $signed(_GEN_28633); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29313 = 6'h6 == state ? $signed(w_15) : $signed(_GEN_28634); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29314 = 6'h6 == state ? $signed(w_16) : $signed(_GEN_28635); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29315 = 6'h6 == state ? $signed(w_17) : $signed(_GEN_28636); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29316 = 6'h6 == state ? $signed(w_18) : $signed(_GEN_28637); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29317 = 6'h6 == state ? $signed(w_19) : $signed(_GEN_28638); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29318 = 6'h6 == state ? $signed(w_20) : $signed(_GEN_28639); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29319 = 6'h6 == state ? $signed(w_21) : $signed(_GEN_28640); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29320 = 6'h6 == state ? $signed(w_22) : $signed(_GEN_28641); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29321 = 6'h6 == state ? $signed(w_23) : $signed(_GEN_28642); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29322 = 6'h6 == state ? $signed(w_24) : $signed(_GEN_28643); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29323 = 6'h6 == state ? $signed(w_25) : $signed(_GEN_28644); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29324 = 6'h6 == state ? $signed(w_26) : $signed(_GEN_28645); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29325 = 6'h6 == state ? $signed(w_27) : $signed(_GEN_28646); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29326 = 6'h6 == state ? $signed(w_28) : $signed(_GEN_28647); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29327 = 6'h6 == state ? $signed(w_29) : $signed(_GEN_28648); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29328 = 6'h6 == state ? $signed(w_30) : $signed(_GEN_28649); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29329 = 6'h6 == state ? $signed(w_31) : $signed(_GEN_28650); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29330 = 6'h6 == state ? $signed(w_32) : $signed(_GEN_28651); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29331 = 6'h6 == state ? $signed(w_33) : $signed(_GEN_28652); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29332 = 6'h6 == state ? $signed(w_34) : $signed(_GEN_28653); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29333 = 6'h6 == state ? $signed(w_35) : $signed(_GEN_28654); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29334 = 6'h6 == state ? $signed(w_36) : $signed(_GEN_28655); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29335 = 6'h6 == state ? $signed(w_37) : $signed(_GEN_28656); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29336 = 6'h6 == state ? $signed(w_38) : $signed(_GEN_28657); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29337 = 6'h6 == state ? $signed(w_39) : $signed(_GEN_28658); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29338 = 6'h6 == state ? $signed(w_40) : $signed(_GEN_28659); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29339 = 6'h6 == state ? $signed(w_41) : $signed(_GEN_28660); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29340 = 6'h6 == state ? $signed(w_42) : $signed(_GEN_28661); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29341 = 6'h6 == state ? $signed(w_43) : $signed(_GEN_28662); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29342 = 6'h6 == state ? $signed(w_44) : $signed(_GEN_28663); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29343 = 6'h6 == state ? $signed(w_45) : $signed(_GEN_28664); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29344 = 6'h6 == state ? $signed(w_46) : $signed(_GEN_28665); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29345 = 6'h6 == state ? $signed(w_47) : $signed(_GEN_28666); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29346 = 6'h6 == state ? $signed(w_48) : $signed(_GEN_28667); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29347 = 6'h6 == state ? $signed(w_49) : $signed(_GEN_28668); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29348 = 6'h6 == state ? $signed(w_50) : $signed(_GEN_28669); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29349 = 6'h6 == state ? $signed(w_51) : $signed(_GEN_28670); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29350 = 6'h6 == state ? $signed(w_52) : $signed(_GEN_28671); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29351 = 6'h6 == state ? $signed(w_53) : $signed(_GEN_28672); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29352 = 6'h6 == state ? $signed(w_54) : $signed(_GEN_28673); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29353 = 6'h6 == state ? $signed(w_55) : $signed(_GEN_28674); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29354 = 6'h6 == state ? $signed(w_56) : $signed(_GEN_28675); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29355 = 6'h6 == state ? $signed(w_57) : $signed(_GEN_28676); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29356 = 6'h6 == state ? $signed(w_58) : $signed(_GEN_28677); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29357 = 6'h6 == state ? $signed(w_59) : $signed(_GEN_28678); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29358 = 6'h6 == state ? $signed(w_60) : $signed(_GEN_28679); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29359 = 6'h6 == state ? $signed(w_61) : $signed(_GEN_28680); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29360 = 6'h6 == state ? $signed(w_62) : $signed(_GEN_28681); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29361 = 6'h6 == state ? $signed(w_63) : $signed(_GEN_28682); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29362 = 6'h6 == state ? $signed(w_64) : $signed(_GEN_28683); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29363 = 6'h6 == state ? $signed(w_65) : $signed(_GEN_28684); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29364 = 6'h6 == state ? $signed(w_66) : $signed(_GEN_28685); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29365 = 6'h6 == state ? $signed(w_67) : $signed(_GEN_28686); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29366 = 6'h6 == state ? $signed(w_68) : $signed(_GEN_28687); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29367 = 6'h6 == state ? $signed(w_69) : $signed(_GEN_28688); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29368 = 6'h6 == state ? $signed(w_70) : $signed(_GEN_28689); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29369 = 6'h6 == state ? $signed(w_71) : $signed(_GEN_28690); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29370 = 6'h6 == state ? $signed(w_72) : $signed(_GEN_28691); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29371 = 6'h6 == state ? $signed(w_73) : $signed(_GEN_28692); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29372 = 6'h6 == state ? $signed(w_74) : $signed(_GEN_28693); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29373 = 6'h6 == state ? $signed(w_75) : $signed(_GEN_28694); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29374 = 6'h6 == state ? $signed(w_76) : $signed(_GEN_28695); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29375 = 6'h6 == state ? $signed(w_77) : $signed(_GEN_28696); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29376 = 6'h6 == state ? $signed(w_78) : $signed(_GEN_28697); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29377 = 6'h6 == state ? $signed(w_79) : $signed(_GEN_28698); // @[digest.scala 40:16 81:19]
  wire  _GEN_29378 = 6'h6 == state ? 1'h0 : _GEN_28699; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_29381 = 6'h6 == state ? $signed(t) : $signed(_GEN_28702); // @[digest.scala 35:16 81:19]
  wire  _GEN_29382 = 6'h6 == state ? 1'h0 : _GEN_28703; // @[digest.scala 81:19 48:24]
  wire  _GEN_29385 = 6'h6 == state ? 1'h0 : _GEN_28706; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_29469 = 6'h6 == state ? $signed(digest_0) : $signed(_GEN_28790); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29470 = 6'h6 == state ? $signed(digest_1) : $signed(_GEN_28791); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29471 = 6'h6 == state ? $signed(digest_2) : $signed(_GEN_28792); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29472 = 6'h6 == state ? $signed(digest_3) : $signed(_GEN_28793); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29473 = 6'h6 == state ? $signed(digest_4) : $signed(_GEN_28794); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29474 = 6'h6 == state ? $signed(digest_5) : $signed(_GEN_28795); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29475 = 6'h6 == state ? $signed(digest_6) : $signed(_GEN_28796); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29476 = 6'h6 == state ? $signed(digest_7) : $signed(_GEN_28797); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29477 = 6'h6 == state ? $signed(digest_8) : $signed(_GEN_28798); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29478 = 6'h6 == state ? $signed(digest_9) : $signed(_GEN_28799); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29479 = 6'h6 == state ? $signed(digest_10) : $signed(_GEN_28800); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29480 = 6'h6 == state ? $signed(digest_11) : $signed(_GEN_28801); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29481 = 6'h6 == state ? $signed(digest_12) : $signed(_GEN_28802); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29482 = 6'h6 == state ? $signed(digest_13) : $signed(_GEN_28803); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29483 = 6'h6 == state ? $signed(digest_14) : $signed(_GEN_28804); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29484 = 6'h6 == state ? $signed(digest_15) : $signed(_GEN_28805); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29485 = 6'h6 == state ? $signed(digest_16) : $signed(_GEN_28806); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29486 = 6'h6 == state ? $signed(digest_17) : $signed(_GEN_28807); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29487 = 6'h6 == state ? $signed(digest_18) : $signed(_GEN_28808); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29488 = 6'h6 == state ? $signed(digest_19) : $signed(_GEN_28809); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29489 = 6'h6 == state ? $signed(digest_20) : $signed(_GEN_28810); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29490 = 6'h6 == state ? $signed(digest_21) : $signed(_GEN_28811); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29491 = 6'h6 == state ? $signed(digest_22) : $signed(_GEN_28812); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29492 = 6'h6 == state ? $signed(digest_23) : $signed(_GEN_28813); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29493 = 6'h6 == state ? $signed(digest_24) : $signed(_GEN_28814); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29494 = 6'h6 == state ? $signed(digest_25) : $signed(_GEN_28815); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29495 = 6'h6 == state ? $signed(digest_26) : $signed(_GEN_28816); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29496 = 6'h6 == state ? $signed(digest_27) : $signed(_GEN_28817); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29497 = 6'h6 == state ? $signed(digest_28) : $signed(_GEN_28818); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29498 = 6'h6 == state ? $signed(digest_29) : $signed(_GEN_28819); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29499 = 6'h6 == state ? $signed(digest_30) : $signed(_GEN_28820); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29500 = 6'h6 == state ? $signed(digest_31) : $signed(_GEN_28821); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29501 = 6'h6 == state ? $signed(digest_32) : $signed(_GEN_28822); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29502 = 6'h6 == state ? $signed(digest_33) : $signed(_GEN_28823); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29503 = 6'h6 == state ? $signed(digest_34) : $signed(_GEN_28824); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29504 = 6'h6 == state ? $signed(digest_35) : $signed(_GEN_28825); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29505 = 6'h6 == state ? $signed(digest_36) : $signed(_GEN_28826); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29506 = 6'h6 == state ? $signed(digest_37) : $signed(_GEN_28827); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29507 = 6'h6 == state ? $signed(digest_38) : $signed(_GEN_28828); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29508 = 6'h6 == state ? $signed(digest_39) : $signed(_GEN_28829); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29509 = 6'h6 == state ? $signed(digest_40) : $signed(_GEN_28830); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29510 = 6'h6 == state ? $signed(digest_41) : $signed(_GEN_28831); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29511 = 6'h6 == state ? $signed(digest_42) : $signed(_GEN_28832); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29512 = 6'h6 == state ? $signed(digest_43) : $signed(_GEN_28833); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29513 = 6'h6 == state ? $signed(digest_44) : $signed(_GEN_28834); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29514 = 6'h6 == state ? $signed(digest_45) : $signed(_GEN_28835); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29515 = 6'h6 == state ? $signed(digest_46) : $signed(_GEN_28836); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29516 = 6'h6 == state ? $signed(digest_47) : $signed(_GEN_28837); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29517 = 6'h6 == state ? $signed(digest_48) : $signed(_GEN_28838); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29518 = 6'h6 == state ? $signed(digest_49) : $signed(_GEN_28839); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29519 = 6'h6 == state ? $signed(digest_50) : $signed(_GEN_28840); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29520 = 6'h6 == state ? $signed(digest_51) : $signed(_GEN_28841); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29521 = 6'h6 == state ? $signed(digest_52) : $signed(_GEN_28842); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29522 = 6'h6 == state ? $signed(digest_53) : $signed(_GEN_28843); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29523 = 6'h6 == state ? $signed(digest_54) : $signed(_GEN_28844); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29524 = 6'h6 == state ? $signed(digest_55) : $signed(_GEN_28845); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29525 = 6'h6 == state ? $signed(digest_56) : $signed(_GEN_28846); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29526 = 6'h6 == state ? $signed(digest_57) : $signed(_GEN_28847); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29527 = 6'h6 == state ? $signed(digest_58) : $signed(_GEN_28848); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29528 = 6'h6 == state ? $signed(digest_59) : $signed(_GEN_28849); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29529 = 6'h6 == state ? $signed(digest_60) : $signed(_GEN_28850); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29530 = 6'h6 == state ? $signed(digest_61) : $signed(_GEN_28851); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29531 = 6'h6 == state ? $signed(digest_62) : $signed(_GEN_28852); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29532 = 6'h6 == state ? $signed(digest_63) : $signed(_GEN_28853); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29533 = 6'h6 == state ? $signed(digest_64) : $signed(_GEN_28854); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29534 = 6'h6 == state ? $signed(digest_65) : $signed(_GEN_28855); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29535 = 6'h6 == state ? $signed(digest_66) : $signed(_GEN_28856); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29536 = 6'h6 == state ? $signed(digest_67) : $signed(_GEN_28857); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29537 = 6'h6 == state ? $signed(digest_68) : $signed(_GEN_28858); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29538 = 6'h6 == state ? $signed(digest_69) : $signed(_GEN_28859); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29539 = 6'h6 == state ? $signed(digest_70) : $signed(_GEN_28860); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29540 = 6'h6 == state ? $signed(digest_71) : $signed(_GEN_28861); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29541 = 6'h6 == state ? $signed(digest_72) : $signed(_GEN_28862); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29542 = 6'h6 == state ? $signed(digest_73) : $signed(_GEN_28863); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29543 = 6'h6 == state ? $signed(digest_74) : $signed(_GEN_28864); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29544 = 6'h6 == state ? $signed(digest_75) : $signed(_GEN_28865); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29545 = 6'h6 == state ? $signed(digest_76) : $signed(_GEN_28866); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29546 = 6'h6 == state ? $signed(digest_77) : $signed(_GEN_28867); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29547 = 6'h6 == state ? $signed(digest_78) : $signed(_GEN_28868); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_29548 = 6'h6 == state ? $signed(digest_79) : $signed(_GEN_28869); // @[digest.scala 81:19 53:21]
  wire  _GEN_29550 = 6'h6 == state ? 1'h0 : _GEN_28871; // @[digest.scala 81:19 58:25]
  wire  _GEN_29633 = 6'h6 == state ? 1'h0 : _GEN_28954; // @[digest.scala 81:19 63:25]
  wire  _GEN_29716 = 6'h6 == state ? 1'h0 : _GEN_29037; // @[digest.scala 81:19 68:25]
  wire  _GEN_29799 = 6'h6 == state ? 1'h0 : _GEN_29120; // @[digest.scala 81:19 73:25]
  wire  _GEN_29882 = 6'h6 == state ? 1'h0 : _GEN_29203; // @[digest.scala 81:19 78:25]
  wire [31:0] _GEN_29883 = 6'h5 == state ? $signed(_GEN_241) : $signed(_GEN_29207); // @[digest.scala 81:19]
  wire [31:0] _GEN_29884 = 6'h5 == state ? $signed(_GEN_242) : $signed(_GEN_29208); // @[digest.scala 81:19]
  wire [31:0] _GEN_29885 = 6'h5 == state ? $signed(_GEN_243) : $signed(_GEN_29209); // @[digest.scala 81:19]
  wire [31:0] _GEN_29886 = 6'h5 == state ? $signed(_GEN_244) : $signed(_GEN_29210); // @[digest.scala 81:19]
  wire [31:0] _GEN_29887 = 6'h5 == state ? $signed(_GEN_245) : $signed(_GEN_29211); // @[digest.scala 81:19]
  wire [31:0] _GEN_29888 = 6'h5 == state ? $signed(_GEN_246) : $signed(_GEN_29212); // @[digest.scala 81:19]
  wire [31:0] _GEN_29889 = 6'h5 == state ? $signed(_GEN_247) : $signed(_GEN_29213); // @[digest.scala 81:19]
  wire [31:0] _GEN_29890 = 6'h5 == state ? $signed(_GEN_248) : $signed(_GEN_29214); // @[digest.scala 81:19]
  wire [31:0] _GEN_29891 = 6'h5 == state ? $signed(_GEN_249) : $signed(_GEN_29215); // @[digest.scala 81:19]
  wire [31:0] _GEN_29892 = 6'h5 == state ? $signed(_GEN_250) : $signed(_GEN_29216); // @[digest.scala 81:19]
  wire [31:0] _GEN_29893 = 6'h5 == state ? $signed(_GEN_251) : $signed(_GEN_29217); // @[digest.scala 81:19]
  wire [31:0] _GEN_29894 = 6'h5 == state ? $signed(_GEN_252) : $signed(_GEN_29218); // @[digest.scala 81:19]
  wire [31:0] _GEN_29895 = 6'h5 == state ? $signed(_GEN_253) : $signed(_GEN_29219); // @[digest.scala 81:19]
  wire [31:0] _GEN_29896 = 6'h5 == state ? $signed(_GEN_254) : $signed(_GEN_29220); // @[digest.scala 81:19]
  wire [31:0] _GEN_29897 = 6'h5 == state ? $signed(_GEN_255) : $signed(_GEN_29221); // @[digest.scala 81:19]
  wire [31:0] _GEN_29898 = 6'h5 == state ? $signed(_GEN_256) : $signed(_GEN_29222); // @[digest.scala 81:19]
  wire [31:0] _GEN_29899 = 6'h5 == state ? $signed(_GEN_257) : $signed(_GEN_29223); // @[digest.scala 81:19]
  wire [31:0] _GEN_29900 = 6'h5 == state ? $signed(_GEN_258) : $signed(_GEN_29224); // @[digest.scala 81:19]
  wire [31:0] _GEN_29901 = 6'h5 == state ? $signed(_GEN_259) : $signed(_GEN_29225); // @[digest.scala 81:19]
  wire [31:0] _GEN_29902 = 6'h5 == state ? $signed(_GEN_260) : $signed(_GEN_29226); // @[digest.scala 81:19]
  wire [31:0] _GEN_29903 = 6'h5 == state ? $signed(_GEN_261) : $signed(_GEN_29227); // @[digest.scala 81:19]
  wire [31:0] _GEN_29904 = 6'h5 == state ? $signed(_GEN_262) : $signed(_GEN_29228); // @[digest.scala 81:19]
  wire [31:0] _GEN_29905 = 6'h5 == state ? $signed(_GEN_263) : $signed(_GEN_29229); // @[digest.scala 81:19]
  wire [31:0] _GEN_29906 = 6'h5 == state ? $signed(_GEN_264) : $signed(_GEN_29230); // @[digest.scala 81:19]
  wire [31:0] _GEN_29907 = 6'h5 == state ? $signed(_GEN_265) : $signed(_GEN_29231); // @[digest.scala 81:19]
  wire [31:0] _GEN_29908 = 6'h5 == state ? $signed(_GEN_266) : $signed(_GEN_29232); // @[digest.scala 81:19]
  wire [31:0] _GEN_29909 = 6'h5 == state ? $signed(_GEN_267) : $signed(_GEN_29233); // @[digest.scala 81:19]
  wire [31:0] _GEN_29910 = 6'h5 == state ? $signed(_GEN_268) : $signed(_GEN_29234); // @[digest.scala 81:19]
  wire [31:0] _GEN_29911 = 6'h5 == state ? $signed(_GEN_269) : $signed(_GEN_29235); // @[digest.scala 81:19]
  wire [31:0] _GEN_29912 = 6'h5 == state ? $signed(_GEN_270) : $signed(_GEN_29236); // @[digest.scala 81:19]
  wire [31:0] _GEN_29913 = 6'h5 == state ? $signed(_GEN_271) : $signed(_GEN_29237); // @[digest.scala 81:19]
  wire [31:0] _GEN_29914 = 6'h5 == state ? $signed(_GEN_272) : $signed(_GEN_29238); // @[digest.scala 81:19]
  wire [31:0] _GEN_29915 = 6'h5 == state ? $signed(_GEN_273) : $signed(_GEN_29239); // @[digest.scala 81:19]
  wire [31:0] _GEN_29916 = 6'h5 == state ? $signed(_GEN_274) : $signed(_GEN_29240); // @[digest.scala 81:19]
  wire [31:0] _GEN_29917 = 6'h5 == state ? $signed(_GEN_275) : $signed(_GEN_29241); // @[digest.scala 81:19]
  wire [31:0] _GEN_29918 = 6'h5 == state ? $signed(_GEN_276) : $signed(_GEN_29242); // @[digest.scala 81:19]
  wire [31:0] _GEN_29919 = 6'h5 == state ? $signed(_GEN_277) : $signed(_GEN_29243); // @[digest.scala 81:19]
  wire [31:0] _GEN_29920 = 6'h5 == state ? $signed(_GEN_278) : $signed(_GEN_29244); // @[digest.scala 81:19]
  wire [31:0] _GEN_29921 = 6'h5 == state ? $signed(_GEN_279) : $signed(_GEN_29245); // @[digest.scala 81:19]
  wire [31:0] _GEN_29922 = 6'h5 == state ? $signed(_GEN_280) : $signed(_GEN_29246); // @[digest.scala 81:19]
  wire [31:0] _GEN_29923 = 6'h5 == state ? $signed(_GEN_281) : $signed(_GEN_29247); // @[digest.scala 81:19]
  wire [31:0] _GEN_29924 = 6'h5 == state ? $signed(_GEN_282) : $signed(_GEN_29248); // @[digest.scala 81:19]
  wire [31:0] _GEN_29925 = 6'h5 == state ? $signed(_GEN_283) : $signed(_GEN_29249); // @[digest.scala 81:19]
  wire [31:0] _GEN_29926 = 6'h5 == state ? $signed(_GEN_284) : $signed(_GEN_29250); // @[digest.scala 81:19]
  wire [31:0] _GEN_29927 = 6'h5 == state ? $signed(_GEN_285) : $signed(_GEN_29251); // @[digest.scala 81:19]
  wire [31:0] _GEN_29928 = 6'h5 == state ? $signed(_GEN_286) : $signed(_GEN_29252); // @[digest.scala 81:19]
  wire [31:0] _GEN_29929 = 6'h5 == state ? $signed(_GEN_287) : $signed(_GEN_29253); // @[digest.scala 81:19]
  wire [31:0] _GEN_29930 = 6'h5 == state ? $signed(_GEN_288) : $signed(_GEN_29254); // @[digest.scala 81:19]
  wire [31:0] _GEN_29931 = 6'h5 == state ? $signed(_GEN_289) : $signed(_GEN_29255); // @[digest.scala 81:19]
  wire [31:0] _GEN_29932 = 6'h5 == state ? $signed(_GEN_290) : $signed(_GEN_29256); // @[digest.scala 81:19]
  wire [31:0] _GEN_29933 = 6'h5 == state ? $signed(_GEN_291) : $signed(_GEN_29257); // @[digest.scala 81:19]
  wire [31:0] _GEN_29934 = 6'h5 == state ? $signed(_GEN_292) : $signed(_GEN_29258); // @[digest.scala 81:19]
  wire [31:0] _GEN_29935 = 6'h5 == state ? $signed(_GEN_293) : $signed(_GEN_29259); // @[digest.scala 81:19]
  wire [31:0] _GEN_29936 = 6'h5 == state ? $signed(_GEN_294) : $signed(_GEN_29260); // @[digest.scala 81:19]
  wire [31:0] _GEN_29937 = 6'h5 == state ? $signed(_GEN_295) : $signed(_GEN_29261); // @[digest.scala 81:19]
  wire [31:0] _GEN_29938 = 6'h5 == state ? $signed(_GEN_296) : $signed(_GEN_29262); // @[digest.scala 81:19]
  wire [31:0] _GEN_29939 = 6'h5 == state ? $signed(_GEN_297) : $signed(_GEN_29263); // @[digest.scala 81:19]
  wire [31:0] _GEN_29940 = 6'h5 == state ? $signed(_GEN_298) : $signed(_GEN_29264); // @[digest.scala 81:19]
  wire [31:0] _GEN_29941 = 6'h5 == state ? $signed(_GEN_299) : $signed(_GEN_29265); // @[digest.scala 81:19]
  wire [31:0] _GEN_29942 = 6'h5 == state ? $signed(_GEN_300) : $signed(_GEN_29266); // @[digest.scala 81:19]
  wire [31:0] _GEN_29943 = 6'h5 == state ? $signed(_GEN_301) : $signed(_GEN_29267); // @[digest.scala 81:19]
  wire [31:0] _GEN_29944 = 6'h5 == state ? $signed(_GEN_302) : $signed(_GEN_29268); // @[digest.scala 81:19]
  wire [31:0] _GEN_29945 = 6'h5 == state ? $signed(_GEN_303) : $signed(_GEN_29269); // @[digest.scala 81:19]
  wire [31:0] _GEN_29946 = 6'h5 == state ? $signed(_GEN_304) : $signed(_GEN_29270); // @[digest.scala 81:19]
  wire [31:0] _GEN_29947 = 6'h5 == state ? $signed(_GEN_305) : $signed(_GEN_29271); // @[digest.scala 81:19]
  wire [31:0] _GEN_29948 = 6'h5 == state ? $signed(_GEN_306) : $signed(_GEN_29272); // @[digest.scala 81:19]
  wire [31:0] _GEN_29949 = 6'h5 == state ? $signed(_GEN_307) : $signed(_GEN_29273); // @[digest.scala 81:19]
  wire [31:0] _GEN_29950 = 6'h5 == state ? $signed(_GEN_308) : $signed(_GEN_29274); // @[digest.scala 81:19]
  wire [31:0] _GEN_29951 = 6'h5 == state ? $signed(_GEN_309) : $signed(_GEN_29275); // @[digest.scala 81:19]
  wire [31:0] _GEN_29952 = 6'h5 == state ? $signed(_GEN_310) : $signed(_GEN_29276); // @[digest.scala 81:19]
  wire [31:0] _GEN_29953 = 6'h5 == state ? $signed(_GEN_311) : $signed(_GEN_29277); // @[digest.scala 81:19]
  wire [31:0] _GEN_29954 = 6'h5 == state ? $signed(_GEN_312) : $signed(_GEN_29278); // @[digest.scala 81:19]
  wire [31:0] _GEN_29955 = 6'h5 == state ? $signed(_GEN_313) : $signed(_GEN_29279); // @[digest.scala 81:19]
  wire [31:0] _GEN_29956 = 6'h5 == state ? $signed(_GEN_314) : $signed(_GEN_29280); // @[digest.scala 81:19]
  wire [31:0] _GEN_29957 = 6'h5 == state ? $signed(_GEN_315) : $signed(_GEN_29281); // @[digest.scala 81:19]
  wire [31:0] _GEN_29958 = 6'h5 == state ? $signed(_GEN_316) : $signed(_GEN_29282); // @[digest.scala 81:19]
  wire [31:0] _GEN_29959 = 6'h5 == state ? $signed(_GEN_317) : $signed(_GEN_29283); // @[digest.scala 81:19]
  wire [31:0] _GEN_29960 = 6'h5 == state ? $signed(_GEN_318) : $signed(_GEN_29284); // @[digest.scala 81:19]
  wire [31:0] _GEN_29961 = 6'h5 == state ? $signed(_GEN_319) : $signed(_GEN_29285); // @[digest.scala 81:19]
  wire [31:0] _GEN_29962 = 6'h5 == state ? $signed(_GEN_320) : $signed(_GEN_29286); // @[digest.scala 81:19]
  wire [5:0] _GEN_29963 = 6'h5 == state ? 6'h6 : _GEN_29205; // @[digest.scala 106:19 81:19]
  wire [31:0] _GEN_29964 = 6'h5 == state ? $signed(i) : $signed(_GEN_29204); // @[digest.scala 23:16 81:19]
  wire [62:0] _GEN_29965 = 6'h5 == state ? $signed({{31{temp[31]}},temp}) : $signed(_GEN_29206); // @[digest.scala 38:19 81:19]
  wire [31:0] _GEN_29966 = 6'h5 == state ? $signed(a) : $signed(_GEN_29287); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_29967 = 6'h5 == state ? $signed(b) : $signed(_GEN_29288); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_29968 = 6'h5 == state ? $signed(c) : $signed(_GEN_29289); // @[digest.scala 26:16 81:19]
  wire [31:0] _GEN_29969 = 6'h5 == state ? $signed(d) : $signed(_GEN_29290); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_29970 = 6'h5 == state ? $signed(e) : $signed(_GEN_29291); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_29971 = 6'h5 == state ? $signed(olda) : $signed(_GEN_29292); // @[digest.scala 29:19 81:19]
  wire [31:0] _GEN_29972 = 6'h5 == state ? $signed(oldb) : $signed(_GEN_29293); // @[digest.scala 30:19 81:19]
  wire [31:0] _GEN_29973 = 6'h5 == state ? $signed(oldc) : $signed(_GEN_29294); // @[digest.scala 31:19 81:19]
  wire [31:0] _GEN_29974 = 6'h5 == state ? $signed(oldd) : $signed(_GEN_29295); // @[digest.scala 32:19 81:19]
  wire [31:0] _GEN_29975 = 6'h5 == state ? $signed(olde) : $signed(_GEN_29296); // @[digest.scala 33:19 81:19]
  wire [31:0] _GEN_29976 = 6'h5 == state ? $signed(j) : $signed(_GEN_29297); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_29977 = 6'h5 == state ? $signed(w_0) : $signed(_GEN_29298); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29978 = 6'h5 == state ? $signed(w_1) : $signed(_GEN_29299); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29979 = 6'h5 == state ? $signed(w_2) : $signed(_GEN_29300); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29980 = 6'h5 == state ? $signed(w_3) : $signed(_GEN_29301); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29981 = 6'h5 == state ? $signed(w_4) : $signed(_GEN_29302); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29982 = 6'h5 == state ? $signed(w_5) : $signed(_GEN_29303); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29983 = 6'h5 == state ? $signed(w_6) : $signed(_GEN_29304); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29984 = 6'h5 == state ? $signed(w_7) : $signed(_GEN_29305); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29985 = 6'h5 == state ? $signed(w_8) : $signed(_GEN_29306); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29986 = 6'h5 == state ? $signed(w_9) : $signed(_GEN_29307); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29987 = 6'h5 == state ? $signed(w_10) : $signed(_GEN_29308); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29988 = 6'h5 == state ? $signed(w_11) : $signed(_GEN_29309); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29989 = 6'h5 == state ? $signed(w_12) : $signed(_GEN_29310); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29990 = 6'h5 == state ? $signed(w_13) : $signed(_GEN_29311); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29991 = 6'h5 == state ? $signed(w_14) : $signed(_GEN_29312); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29992 = 6'h5 == state ? $signed(w_15) : $signed(_GEN_29313); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29993 = 6'h5 == state ? $signed(w_16) : $signed(_GEN_29314); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29994 = 6'h5 == state ? $signed(w_17) : $signed(_GEN_29315); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29995 = 6'h5 == state ? $signed(w_18) : $signed(_GEN_29316); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29996 = 6'h5 == state ? $signed(w_19) : $signed(_GEN_29317); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29997 = 6'h5 == state ? $signed(w_20) : $signed(_GEN_29318); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29998 = 6'h5 == state ? $signed(w_21) : $signed(_GEN_29319); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_29999 = 6'h5 == state ? $signed(w_22) : $signed(_GEN_29320); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30000 = 6'h5 == state ? $signed(w_23) : $signed(_GEN_29321); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30001 = 6'h5 == state ? $signed(w_24) : $signed(_GEN_29322); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30002 = 6'h5 == state ? $signed(w_25) : $signed(_GEN_29323); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30003 = 6'h5 == state ? $signed(w_26) : $signed(_GEN_29324); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30004 = 6'h5 == state ? $signed(w_27) : $signed(_GEN_29325); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30005 = 6'h5 == state ? $signed(w_28) : $signed(_GEN_29326); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30006 = 6'h5 == state ? $signed(w_29) : $signed(_GEN_29327); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30007 = 6'h5 == state ? $signed(w_30) : $signed(_GEN_29328); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30008 = 6'h5 == state ? $signed(w_31) : $signed(_GEN_29329); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30009 = 6'h5 == state ? $signed(w_32) : $signed(_GEN_29330); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30010 = 6'h5 == state ? $signed(w_33) : $signed(_GEN_29331); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30011 = 6'h5 == state ? $signed(w_34) : $signed(_GEN_29332); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30012 = 6'h5 == state ? $signed(w_35) : $signed(_GEN_29333); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30013 = 6'h5 == state ? $signed(w_36) : $signed(_GEN_29334); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30014 = 6'h5 == state ? $signed(w_37) : $signed(_GEN_29335); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30015 = 6'h5 == state ? $signed(w_38) : $signed(_GEN_29336); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30016 = 6'h5 == state ? $signed(w_39) : $signed(_GEN_29337); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30017 = 6'h5 == state ? $signed(w_40) : $signed(_GEN_29338); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30018 = 6'h5 == state ? $signed(w_41) : $signed(_GEN_29339); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30019 = 6'h5 == state ? $signed(w_42) : $signed(_GEN_29340); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30020 = 6'h5 == state ? $signed(w_43) : $signed(_GEN_29341); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30021 = 6'h5 == state ? $signed(w_44) : $signed(_GEN_29342); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30022 = 6'h5 == state ? $signed(w_45) : $signed(_GEN_29343); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30023 = 6'h5 == state ? $signed(w_46) : $signed(_GEN_29344); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30024 = 6'h5 == state ? $signed(w_47) : $signed(_GEN_29345); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30025 = 6'h5 == state ? $signed(w_48) : $signed(_GEN_29346); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30026 = 6'h5 == state ? $signed(w_49) : $signed(_GEN_29347); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30027 = 6'h5 == state ? $signed(w_50) : $signed(_GEN_29348); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30028 = 6'h5 == state ? $signed(w_51) : $signed(_GEN_29349); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30029 = 6'h5 == state ? $signed(w_52) : $signed(_GEN_29350); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30030 = 6'h5 == state ? $signed(w_53) : $signed(_GEN_29351); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30031 = 6'h5 == state ? $signed(w_54) : $signed(_GEN_29352); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30032 = 6'h5 == state ? $signed(w_55) : $signed(_GEN_29353); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30033 = 6'h5 == state ? $signed(w_56) : $signed(_GEN_29354); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30034 = 6'h5 == state ? $signed(w_57) : $signed(_GEN_29355); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30035 = 6'h5 == state ? $signed(w_58) : $signed(_GEN_29356); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30036 = 6'h5 == state ? $signed(w_59) : $signed(_GEN_29357); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30037 = 6'h5 == state ? $signed(w_60) : $signed(_GEN_29358); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30038 = 6'h5 == state ? $signed(w_61) : $signed(_GEN_29359); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30039 = 6'h5 == state ? $signed(w_62) : $signed(_GEN_29360); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30040 = 6'h5 == state ? $signed(w_63) : $signed(_GEN_29361); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30041 = 6'h5 == state ? $signed(w_64) : $signed(_GEN_29362); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30042 = 6'h5 == state ? $signed(w_65) : $signed(_GEN_29363); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30043 = 6'h5 == state ? $signed(w_66) : $signed(_GEN_29364); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30044 = 6'h5 == state ? $signed(w_67) : $signed(_GEN_29365); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30045 = 6'h5 == state ? $signed(w_68) : $signed(_GEN_29366); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30046 = 6'h5 == state ? $signed(w_69) : $signed(_GEN_29367); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30047 = 6'h5 == state ? $signed(w_70) : $signed(_GEN_29368); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30048 = 6'h5 == state ? $signed(w_71) : $signed(_GEN_29369); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30049 = 6'h5 == state ? $signed(w_72) : $signed(_GEN_29370); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30050 = 6'h5 == state ? $signed(w_73) : $signed(_GEN_29371); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30051 = 6'h5 == state ? $signed(w_74) : $signed(_GEN_29372); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30052 = 6'h5 == state ? $signed(w_75) : $signed(_GEN_29373); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30053 = 6'h5 == state ? $signed(w_76) : $signed(_GEN_29374); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30054 = 6'h5 == state ? $signed(w_77) : $signed(_GEN_29375); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30055 = 6'h5 == state ? $signed(w_78) : $signed(_GEN_29376); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30056 = 6'h5 == state ? $signed(w_79) : $signed(_GEN_29377); // @[digest.scala 40:16 81:19]
  wire  _GEN_30057 = 6'h5 == state ? 1'h0 : _GEN_29378; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_30060 = 6'h5 == state ? $signed(t) : $signed(_GEN_29381); // @[digest.scala 35:16 81:19]
  wire  _GEN_30061 = 6'h5 == state ? 1'h0 : _GEN_29382; // @[digest.scala 81:19 48:24]
  wire  _GEN_30064 = 6'h5 == state ? 1'h0 : _GEN_29385; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_30148 = 6'h5 == state ? $signed(digest_0) : $signed(_GEN_29469); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30149 = 6'h5 == state ? $signed(digest_1) : $signed(_GEN_29470); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30150 = 6'h5 == state ? $signed(digest_2) : $signed(_GEN_29471); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30151 = 6'h5 == state ? $signed(digest_3) : $signed(_GEN_29472); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30152 = 6'h5 == state ? $signed(digest_4) : $signed(_GEN_29473); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30153 = 6'h5 == state ? $signed(digest_5) : $signed(_GEN_29474); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30154 = 6'h5 == state ? $signed(digest_6) : $signed(_GEN_29475); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30155 = 6'h5 == state ? $signed(digest_7) : $signed(_GEN_29476); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30156 = 6'h5 == state ? $signed(digest_8) : $signed(_GEN_29477); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30157 = 6'h5 == state ? $signed(digest_9) : $signed(_GEN_29478); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30158 = 6'h5 == state ? $signed(digest_10) : $signed(_GEN_29479); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30159 = 6'h5 == state ? $signed(digest_11) : $signed(_GEN_29480); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30160 = 6'h5 == state ? $signed(digest_12) : $signed(_GEN_29481); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30161 = 6'h5 == state ? $signed(digest_13) : $signed(_GEN_29482); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30162 = 6'h5 == state ? $signed(digest_14) : $signed(_GEN_29483); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30163 = 6'h5 == state ? $signed(digest_15) : $signed(_GEN_29484); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30164 = 6'h5 == state ? $signed(digest_16) : $signed(_GEN_29485); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30165 = 6'h5 == state ? $signed(digest_17) : $signed(_GEN_29486); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30166 = 6'h5 == state ? $signed(digest_18) : $signed(_GEN_29487); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30167 = 6'h5 == state ? $signed(digest_19) : $signed(_GEN_29488); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30168 = 6'h5 == state ? $signed(digest_20) : $signed(_GEN_29489); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30169 = 6'h5 == state ? $signed(digest_21) : $signed(_GEN_29490); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30170 = 6'h5 == state ? $signed(digest_22) : $signed(_GEN_29491); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30171 = 6'h5 == state ? $signed(digest_23) : $signed(_GEN_29492); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30172 = 6'h5 == state ? $signed(digest_24) : $signed(_GEN_29493); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30173 = 6'h5 == state ? $signed(digest_25) : $signed(_GEN_29494); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30174 = 6'h5 == state ? $signed(digest_26) : $signed(_GEN_29495); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30175 = 6'h5 == state ? $signed(digest_27) : $signed(_GEN_29496); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30176 = 6'h5 == state ? $signed(digest_28) : $signed(_GEN_29497); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30177 = 6'h5 == state ? $signed(digest_29) : $signed(_GEN_29498); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30178 = 6'h5 == state ? $signed(digest_30) : $signed(_GEN_29499); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30179 = 6'h5 == state ? $signed(digest_31) : $signed(_GEN_29500); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30180 = 6'h5 == state ? $signed(digest_32) : $signed(_GEN_29501); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30181 = 6'h5 == state ? $signed(digest_33) : $signed(_GEN_29502); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30182 = 6'h5 == state ? $signed(digest_34) : $signed(_GEN_29503); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30183 = 6'h5 == state ? $signed(digest_35) : $signed(_GEN_29504); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30184 = 6'h5 == state ? $signed(digest_36) : $signed(_GEN_29505); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30185 = 6'h5 == state ? $signed(digest_37) : $signed(_GEN_29506); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30186 = 6'h5 == state ? $signed(digest_38) : $signed(_GEN_29507); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30187 = 6'h5 == state ? $signed(digest_39) : $signed(_GEN_29508); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30188 = 6'h5 == state ? $signed(digest_40) : $signed(_GEN_29509); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30189 = 6'h5 == state ? $signed(digest_41) : $signed(_GEN_29510); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30190 = 6'h5 == state ? $signed(digest_42) : $signed(_GEN_29511); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30191 = 6'h5 == state ? $signed(digest_43) : $signed(_GEN_29512); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30192 = 6'h5 == state ? $signed(digest_44) : $signed(_GEN_29513); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30193 = 6'h5 == state ? $signed(digest_45) : $signed(_GEN_29514); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30194 = 6'h5 == state ? $signed(digest_46) : $signed(_GEN_29515); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30195 = 6'h5 == state ? $signed(digest_47) : $signed(_GEN_29516); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30196 = 6'h5 == state ? $signed(digest_48) : $signed(_GEN_29517); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30197 = 6'h5 == state ? $signed(digest_49) : $signed(_GEN_29518); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30198 = 6'h5 == state ? $signed(digest_50) : $signed(_GEN_29519); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30199 = 6'h5 == state ? $signed(digest_51) : $signed(_GEN_29520); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30200 = 6'h5 == state ? $signed(digest_52) : $signed(_GEN_29521); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30201 = 6'h5 == state ? $signed(digest_53) : $signed(_GEN_29522); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30202 = 6'h5 == state ? $signed(digest_54) : $signed(_GEN_29523); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30203 = 6'h5 == state ? $signed(digest_55) : $signed(_GEN_29524); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30204 = 6'h5 == state ? $signed(digest_56) : $signed(_GEN_29525); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30205 = 6'h5 == state ? $signed(digest_57) : $signed(_GEN_29526); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30206 = 6'h5 == state ? $signed(digest_58) : $signed(_GEN_29527); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30207 = 6'h5 == state ? $signed(digest_59) : $signed(_GEN_29528); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30208 = 6'h5 == state ? $signed(digest_60) : $signed(_GEN_29529); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30209 = 6'h5 == state ? $signed(digest_61) : $signed(_GEN_29530); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30210 = 6'h5 == state ? $signed(digest_62) : $signed(_GEN_29531); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30211 = 6'h5 == state ? $signed(digest_63) : $signed(_GEN_29532); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30212 = 6'h5 == state ? $signed(digest_64) : $signed(_GEN_29533); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30213 = 6'h5 == state ? $signed(digest_65) : $signed(_GEN_29534); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30214 = 6'h5 == state ? $signed(digest_66) : $signed(_GEN_29535); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30215 = 6'h5 == state ? $signed(digest_67) : $signed(_GEN_29536); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30216 = 6'h5 == state ? $signed(digest_68) : $signed(_GEN_29537); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30217 = 6'h5 == state ? $signed(digest_69) : $signed(_GEN_29538); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30218 = 6'h5 == state ? $signed(digest_70) : $signed(_GEN_29539); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30219 = 6'h5 == state ? $signed(digest_71) : $signed(_GEN_29540); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30220 = 6'h5 == state ? $signed(digest_72) : $signed(_GEN_29541); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30221 = 6'h5 == state ? $signed(digest_73) : $signed(_GEN_29542); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30222 = 6'h5 == state ? $signed(digest_74) : $signed(_GEN_29543); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30223 = 6'h5 == state ? $signed(digest_75) : $signed(_GEN_29544); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30224 = 6'h5 == state ? $signed(digest_76) : $signed(_GEN_29545); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30225 = 6'h5 == state ? $signed(digest_77) : $signed(_GEN_29546); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30226 = 6'h5 == state ? $signed(digest_78) : $signed(_GEN_29547); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30227 = 6'h5 == state ? $signed(digest_79) : $signed(_GEN_29548); // @[digest.scala 81:19 53:21]
  wire  _GEN_30229 = 6'h5 == state ? 1'h0 : _GEN_29550; // @[digest.scala 81:19 58:25]
  wire  _GEN_30312 = 6'h5 == state ? 1'h0 : _GEN_29633; // @[digest.scala 81:19 63:25]
  wire  _GEN_30395 = 6'h5 == state ? 1'h0 : _GEN_29716; // @[digest.scala 81:19 68:25]
  wire  _GEN_30478 = 6'h5 == state ? 1'h0 : _GEN_29799; // @[digest.scala 81:19 73:25]
  wire  _GEN_30561 = 6'h5 == state ? 1'h0 : _GEN_29882; // @[digest.scala 81:19 78:25]
  wire [62:0] _GEN_30562 = 6'h4 == state ? $signed(_temp_T_9) : $signed(_GEN_29965); // @[digest.scala 101:18 81:19]
  wire [5:0] _GEN_30563 = 6'h4 == state ? 6'h5 : _GEN_29963; // @[digest.scala 102:19 81:19]
  wire [31:0] _GEN_30564 = 6'h4 == state ? $signed(blks_0) : $signed(_GEN_29883); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30565 = 6'h4 == state ? $signed(blks_1) : $signed(_GEN_29884); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30566 = 6'h4 == state ? $signed(blks_2) : $signed(_GEN_29885); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30567 = 6'h4 == state ? $signed(blks_3) : $signed(_GEN_29886); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30568 = 6'h4 == state ? $signed(blks_4) : $signed(_GEN_29887); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30569 = 6'h4 == state ? $signed(blks_5) : $signed(_GEN_29888); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30570 = 6'h4 == state ? $signed(blks_6) : $signed(_GEN_29889); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30571 = 6'h4 == state ? $signed(blks_7) : $signed(_GEN_29890); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30572 = 6'h4 == state ? $signed(blks_8) : $signed(_GEN_29891); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30573 = 6'h4 == state ? $signed(blks_9) : $signed(_GEN_29892); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30574 = 6'h4 == state ? $signed(blks_10) : $signed(_GEN_29893); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30575 = 6'h4 == state ? $signed(blks_11) : $signed(_GEN_29894); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30576 = 6'h4 == state ? $signed(blks_12) : $signed(_GEN_29895); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30577 = 6'h4 == state ? $signed(blks_13) : $signed(_GEN_29896); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30578 = 6'h4 == state ? $signed(blks_14) : $signed(_GEN_29897); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30579 = 6'h4 == state ? $signed(blks_15) : $signed(_GEN_29898); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30580 = 6'h4 == state ? $signed(blks_16) : $signed(_GEN_29899); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30581 = 6'h4 == state ? $signed(blks_17) : $signed(_GEN_29900); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30582 = 6'h4 == state ? $signed(blks_18) : $signed(_GEN_29901); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30583 = 6'h4 == state ? $signed(blks_19) : $signed(_GEN_29902); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30584 = 6'h4 == state ? $signed(blks_20) : $signed(_GEN_29903); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30585 = 6'h4 == state ? $signed(blks_21) : $signed(_GEN_29904); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30586 = 6'h4 == state ? $signed(blks_22) : $signed(_GEN_29905); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30587 = 6'h4 == state ? $signed(blks_23) : $signed(_GEN_29906); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30588 = 6'h4 == state ? $signed(blks_24) : $signed(_GEN_29907); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30589 = 6'h4 == state ? $signed(blks_25) : $signed(_GEN_29908); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30590 = 6'h4 == state ? $signed(blks_26) : $signed(_GEN_29909); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30591 = 6'h4 == state ? $signed(blks_27) : $signed(_GEN_29910); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30592 = 6'h4 == state ? $signed(blks_28) : $signed(_GEN_29911); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30593 = 6'h4 == state ? $signed(blks_29) : $signed(_GEN_29912); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30594 = 6'h4 == state ? $signed(blks_30) : $signed(_GEN_29913); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30595 = 6'h4 == state ? $signed(blks_31) : $signed(_GEN_29914); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30596 = 6'h4 == state ? $signed(blks_32) : $signed(_GEN_29915); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30597 = 6'h4 == state ? $signed(blks_33) : $signed(_GEN_29916); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30598 = 6'h4 == state ? $signed(blks_34) : $signed(_GEN_29917); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30599 = 6'h4 == state ? $signed(blks_35) : $signed(_GEN_29918); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30600 = 6'h4 == state ? $signed(blks_36) : $signed(_GEN_29919); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30601 = 6'h4 == state ? $signed(blks_37) : $signed(_GEN_29920); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30602 = 6'h4 == state ? $signed(blks_38) : $signed(_GEN_29921); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30603 = 6'h4 == state ? $signed(blks_39) : $signed(_GEN_29922); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30604 = 6'h4 == state ? $signed(blks_40) : $signed(_GEN_29923); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30605 = 6'h4 == state ? $signed(blks_41) : $signed(_GEN_29924); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30606 = 6'h4 == state ? $signed(blks_42) : $signed(_GEN_29925); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30607 = 6'h4 == state ? $signed(blks_43) : $signed(_GEN_29926); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30608 = 6'h4 == state ? $signed(blks_44) : $signed(_GEN_29927); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30609 = 6'h4 == state ? $signed(blks_45) : $signed(_GEN_29928); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30610 = 6'h4 == state ? $signed(blks_46) : $signed(_GEN_29929); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30611 = 6'h4 == state ? $signed(blks_47) : $signed(_GEN_29930); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30612 = 6'h4 == state ? $signed(blks_48) : $signed(_GEN_29931); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30613 = 6'h4 == state ? $signed(blks_49) : $signed(_GEN_29932); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30614 = 6'h4 == state ? $signed(blks_50) : $signed(_GEN_29933); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30615 = 6'h4 == state ? $signed(blks_51) : $signed(_GEN_29934); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30616 = 6'h4 == state ? $signed(blks_52) : $signed(_GEN_29935); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30617 = 6'h4 == state ? $signed(blks_53) : $signed(_GEN_29936); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30618 = 6'h4 == state ? $signed(blks_54) : $signed(_GEN_29937); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30619 = 6'h4 == state ? $signed(blks_55) : $signed(_GEN_29938); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30620 = 6'h4 == state ? $signed(blks_56) : $signed(_GEN_29939); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30621 = 6'h4 == state ? $signed(blks_57) : $signed(_GEN_29940); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30622 = 6'h4 == state ? $signed(blks_58) : $signed(_GEN_29941); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30623 = 6'h4 == state ? $signed(blks_59) : $signed(_GEN_29942); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30624 = 6'h4 == state ? $signed(blks_60) : $signed(_GEN_29943); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30625 = 6'h4 == state ? $signed(blks_61) : $signed(_GEN_29944); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30626 = 6'h4 == state ? $signed(blks_62) : $signed(_GEN_29945); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30627 = 6'h4 == state ? $signed(blks_63) : $signed(_GEN_29946); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30628 = 6'h4 == state ? $signed(blks_64) : $signed(_GEN_29947); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30629 = 6'h4 == state ? $signed(blks_65) : $signed(_GEN_29948); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30630 = 6'h4 == state ? $signed(blks_66) : $signed(_GEN_29949); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30631 = 6'h4 == state ? $signed(blks_67) : $signed(_GEN_29950); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30632 = 6'h4 == state ? $signed(blks_68) : $signed(_GEN_29951); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30633 = 6'h4 == state ? $signed(blks_69) : $signed(_GEN_29952); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30634 = 6'h4 == state ? $signed(blks_70) : $signed(_GEN_29953); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30635 = 6'h4 == state ? $signed(blks_71) : $signed(_GEN_29954); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30636 = 6'h4 == state ? $signed(blks_72) : $signed(_GEN_29955); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30637 = 6'h4 == state ? $signed(blks_73) : $signed(_GEN_29956); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30638 = 6'h4 == state ? $signed(blks_74) : $signed(_GEN_29957); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30639 = 6'h4 == state ? $signed(blks_75) : $signed(_GEN_29958); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30640 = 6'h4 == state ? $signed(blks_76) : $signed(_GEN_29959); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30641 = 6'h4 == state ? $signed(blks_77) : $signed(_GEN_29960); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30642 = 6'h4 == state ? $signed(blks_78) : $signed(_GEN_29961); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30643 = 6'h4 == state ? $signed(blks_79) : $signed(_GEN_29962); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_30644 = 6'h4 == state ? $signed(i) : $signed(_GEN_29964); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_30645 = 6'h4 == state ? $signed(a) : $signed(_GEN_29966); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_30646 = 6'h4 == state ? $signed(b) : $signed(_GEN_29967); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_30647 = 6'h4 == state ? $signed(c) : $signed(_GEN_29968); // @[digest.scala 26:16 81:19]
  wire [31:0] _GEN_30648 = 6'h4 == state ? $signed(d) : $signed(_GEN_29969); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_30649 = 6'h4 == state ? $signed(e) : $signed(_GEN_29970); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_30650 = 6'h4 == state ? $signed(olda) : $signed(_GEN_29971); // @[digest.scala 29:19 81:19]
  wire [31:0] _GEN_30651 = 6'h4 == state ? $signed(oldb) : $signed(_GEN_29972); // @[digest.scala 30:19 81:19]
  wire [31:0] _GEN_30652 = 6'h4 == state ? $signed(oldc) : $signed(_GEN_29973); // @[digest.scala 31:19 81:19]
  wire [31:0] _GEN_30653 = 6'h4 == state ? $signed(oldd) : $signed(_GEN_29974); // @[digest.scala 32:19 81:19]
  wire [31:0] _GEN_30654 = 6'h4 == state ? $signed(olde) : $signed(_GEN_29975); // @[digest.scala 33:19 81:19]
  wire [31:0] _GEN_30655 = 6'h4 == state ? $signed(j) : $signed(_GEN_29976); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_30656 = 6'h4 == state ? $signed(w_0) : $signed(_GEN_29977); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30657 = 6'h4 == state ? $signed(w_1) : $signed(_GEN_29978); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30658 = 6'h4 == state ? $signed(w_2) : $signed(_GEN_29979); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30659 = 6'h4 == state ? $signed(w_3) : $signed(_GEN_29980); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30660 = 6'h4 == state ? $signed(w_4) : $signed(_GEN_29981); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30661 = 6'h4 == state ? $signed(w_5) : $signed(_GEN_29982); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30662 = 6'h4 == state ? $signed(w_6) : $signed(_GEN_29983); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30663 = 6'h4 == state ? $signed(w_7) : $signed(_GEN_29984); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30664 = 6'h4 == state ? $signed(w_8) : $signed(_GEN_29985); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30665 = 6'h4 == state ? $signed(w_9) : $signed(_GEN_29986); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30666 = 6'h4 == state ? $signed(w_10) : $signed(_GEN_29987); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30667 = 6'h4 == state ? $signed(w_11) : $signed(_GEN_29988); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30668 = 6'h4 == state ? $signed(w_12) : $signed(_GEN_29989); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30669 = 6'h4 == state ? $signed(w_13) : $signed(_GEN_29990); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30670 = 6'h4 == state ? $signed(w_14) : $signed(_GEN_29991); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30671 = 6'h4 == state ? $signed(w_15) : $signed(_GEN_29992); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30672 = 6'h4 == state ? $signed(w_16) : $signed(_GEN_29993); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30673 = 6'h4 == state ? $signed(w_17) : $signed(_GEN_29994); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30674 = 6'h4 == state ? $signed(w_18) : $signed(_GEN_29995); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30675 = 6'h4 == state ? $signed(w_19) : $signed(_GEN_29996); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30676 = 6'h4 == state ? $signed(w_20) : $signed(_GEN_29997); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30677 = 6'h4 == state ? $signed(w_21) : $signed(_GEN_29998); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30678 = 6'h4 == state ? $signed(w_22) : $signed(_GEN_29999); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30679 = 6'h4 == state ? $signed(w_23) : $signed(_GEN_30000); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30680 = 6'h4 == state ? $signed(w_24) : $signed(_GEN_30001); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30681 = 6'h4 == state ? $signed(w_25) : $signed(_GEN_30002); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30682 = 6'h4 == state ? $signed(w_26) : $signed(_GEN_30003); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30683 = 6'h4 == state ? $signed(w_27) : $signed(_GEN_30004); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30684 = 6'h4 == state ? $signed(w_28) : $signed(_GEN_30005); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30685 = 6'h4 == state ? $signed(w_29) : $signed(_GEN_30006); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30686 = 6'h4 == state ? $signed(w_30) : $signed(_GEN_30007); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30687 = 6'h4 == state ? $signed(w_31) : $signed(_GEN_30008); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30688 = 6'h4 == state ? $signed(w_32) : $signed(_GEN_30009); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30689 = 6'h4 == state ? $signed(w_33) : $signed(_GEN_30010); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30690 = 6'h4 == state ? $signed(w_34) : $signed(_GEN_30011); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30691 = 6'h4 == state ? $signed(w_35) : $signed(_GEN_30012); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30692 = 6'h4 == state ? $signed(w_36) : $signed(_GEN_30013); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30693 = 6'h4 == state ? $signed(w_37) : $signed(_GEN_30014); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30694 = 6'h4 == state ? $signed(w_38) : $signed(_GEN_30015); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30695 = 6'h4 == state ? $signed(w_39) : $signed(_GEN_30016); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30696 = 6'h4 == state ? $signed(w_40) : $signed(_GEN_30017); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30697 = 6'h4 == state ? $signed(w_41) : $signed(_GEN_30018); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30698 = 6'h4 == state ? $signed(w_42) : $signed(_GEN_30019); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30699 = 6'h4 == state ? $signed(w_43) : $signed(_GEN_30020); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30700 = 6'h4 == state ? $signed(w_44) : $signed(_GEN_30021); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30701 = 6'h4 == state ? $signed(w_45) : $signed(_GEN_30022); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30702 = 6'h4 == state ? $signed(w_46) : $signed(_GEN_30023); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30703 = 6'h4 == state ? $signed(w_47) : $signed(_GEN_30024); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30704 = 6'h4 == state ? $signed(w_48) : $signed(_GEN_30025); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30705 = 6'h4 == state ? $signed(w_49) : $signed(_GEN_30026); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30706 = 6'h4 == state ? $signed(w_50) : $signed(_GEN_30027); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30707 = 6'h4 == state ? $signed(w_51) : $signed(_GEN_30028); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30708 = 6'h4 == state ? $signed(w_52) : $signed(_GEN_30029); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30709 = 6'h4 == state ? $signed(w_53) : $signed(_GEN_30030); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30710 = 6'h4 == state ? $signed(w_54) : $signed(_GEN_30031); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30711 = 6'h4 == state ? $signed(w_55) : $signed(_GEN_30032); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30712 = 6'h4 == state ? $signed(w_56) : $signed(_GEN_30033); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30713 = 6'h4 == state ? $signed(w_57) : $signed(_GEN_30034); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30714 = 6'h4 == state ? $signed(w_58) : $signed(_GEN_30035); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30715 = 6'h4 == state ? $signed(w_59) : $signed(_GEN_30036); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30716 = 6'h4 == state ? $signed(w_60) : $signed(_GEN_30037); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30717 = 6'h4 == state ? $signed(w_61) : $signed(_GEN_30038); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30718 = 6'h4 == state ? $signed(w_62) : $signed(_GEN_30039); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30719 = 6'h4 == state ? $signed(w_63) : $signed(_GEN_30040); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30720 = 6'h4 == state ? $signed(w_64) : $signed(_GEN_30041); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30721 = 6'h4 == state ? $signed(w_65) : $signed(_GEN_30042); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30722 = 6'h4 == state ? $signed(w_66) : $signed(_GEN_30043); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30723 = 6'h4 == state ? $signed(w_67) : $signed(_GEN_30044); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30724 = 6'h4 == state ? $signed(w_68) : $signed(_GEN_30045); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30725 = 6'h4 == state ? $signed(w_69) : $signed(_GEN_30046); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30726 = 6'h4 == state ? $signed(w_70) : $signed(_GEN_30047); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30727 = 6'h4 == state ? $signed(w_71) : $signed(_GEN_30048); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30728 = 6'h4 == state ? $signed(w_72) : $signed(_GEN_30049); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30729 = 6'h4 == state ? $signed(w_73) : $signed(_GEN_30050); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30730 = 6'h4 == state ? $signed(w_74) : $signed(_GEN_30051); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30731 = 6'h4 == state ? $signed(w_75) : $signed(_GEN_30052); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30732 = 6'h4 == state ? $signed(w_76) : $signed(_GEN_30053); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30733 = 6'h4 == state ? $signed(w_77) : $signed(_GEN_30054); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30734 = 6'h4 == state ? $signed(w_78) : $signed(_GEN_30055); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_30735 = 6'h4 == state ? $signed(w_79) : $signed(_GEN_30056); // @[digest.scala 40:16 81:19]
  wire  _GEN_30736 = 6'h4 == state ? 1'h0 : _GEN_30057; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_30739 = 6'h4 == state ? $signed(t) : $signed(_GEN_30060); // @[digest.scala 35:16 81:19]
  wire  _GEN_30740 = 6'h4 == state ? 1'h0 : _GEN_30061; // @[digest.scala 81:19 48:24]
  wire  _GEN_30743 = 6'h4 == state ? 1'h0 : _GEN_30064; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_30827 = 6'h4 == state ? $signed(digest_0) : $signed(_GEN_30148); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30828 = 6'h4 == state ? $signed(digest_1) : $signed(_GEN_30149); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30829 = 6'h4 == state ? $signed(digest_2) : $signed(_GEN_30150); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30830 = 6'h4 == state ? $signed(digest_3) : $signed(_GEN_30151); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30831 = 6'h4 == state ? $signed(digest_4) : $signed(_GEN_30152); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30832 = 6'h4 == state ? $signed(digest_5) : $signed(_GEN_30153); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30833 = 6'h4 == state ? $signed(digest_6) : $signed(_GEN_30154); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30834 = 6'h4 == state ? $signed(digest_7) : $signed(_GEN_30155); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30835 = 6'h4 == state ? $signed(digest_8) : $signed(_GEN_30156); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30836 = 6'h4 == state ? $signed(digest_9) : $signed(_GEN_30157); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30837 = 6'h4 == state ? $signed(digest_10) : $signed(_GEN_30158); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30838 = 6'h4 == state ? $signed(digest_11) : $signed(_GEN_30159); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30839 = 6'h4 == state ? $signed(digest_12) : $signed(_GEN_30160); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30840 = 6'h4 == state ? $signed(digest_13) : $signed(_GEN_30161); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30841 = 6'h4 == state ? $signed(digest_14) : $signed(_GEN_30162); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30842 = 6'h4 == state ? $signed(digest_15) : $signed(_GEN_30163); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30843 = 6'h4 == state ? $signed(digest_16) : $signed(_GEN_30164); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30844 = 6'h4 == state ? $signed(digest_17) : $signed(_GEN_30165); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30845 = 6'h4 == state ? $signed(digest_18) : $signed(_GEN_30166); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30846 = 6'h4 == state ? $signed(digest_19) : $signed(_GEN_30167); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30847 = 6'h4 == state ? $signed(digest_20) : $signed(_GEN_30168); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30848 = 6'h4 == state ? $signed(digest_21) : $signed(_GEN_30169); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30849 = 6'h4 == state ? $signed(digest_22) : $signed(_GEN_30170); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30850 = 6'h4 == state ? $signed(digest_23) : $signed(_GEN_30171); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30851 = 6'h4 == state ? $signed(digest_24) : $signed(_GEN_30172); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30852 = 6'h4 == state ? $signed(digest_25) : $signed(_GEN_30173); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30853 = 6'h4 == state ? $signed(digest_26) : $signed(_GEN_30174); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30854 = 6'h4 == state ? $signed(digest_27) : $signed(_GEN_30175); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30855 = 6'h4 == state ? $signed(digest_28) : $signed(_GEN_30176); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30856 = 6'h4 == state ? $signed(digest_29) : $signed(_GEN_30177); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30857 = 6'h4 == state ? $signed(digest_30) : $signed(_GEN_30178); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30858 = 6'h4 == state ? $signed(digest_31) : $signed(_GEN_30179); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30859 = 6'h4 == state ? $signed(digest_32) : $signed(_GEN_30180); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30860 = 6'h4 == state ? $signed(digest_33) : $signed(_GEN_30181); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30861 = 6'h4 == state ? $signed(digest_34) : $signed(_GEN_30182); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30862 = 6'h4 == state ? $signed(digest_35) : $signed(_GEN_30183); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30863 = 6'h4 == state ? $signed(digest_36) : $signed(_GEN_30184); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30864 = 6'h4 == state ? $signed(digest_37) : $signed(_GEN_30185); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30865 = 6'h4 == state ? $signed(digest_38) : $signed(_GEN_30186); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30866 = 6'h4 == state ? $signed(digest_39) : $signed(_GEN_30187); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30867 = 6'h4 == state ? $signed(digest_40) : $signed(_GEN_30188); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30868 = 6'h4 == state ? $signed(digest_41) : $signed(_GEN_30189); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30869 = 6'h4 == state ? $signed(digest_42) : $signed(_GEN_30190); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30870 = 6'h4 == state ? $signed(digest_43) : $signed(_GEN_30191); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30871 = 6'h4 == state ? $signed(digest_44) : $signed(_GEN_30192); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30872 = 6'h4 == state ? $signed(digest_45) : $signed(_GEN_30193); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30873 = 6'h4 == state ? $signed(digest_46) : $signed(_GEN_30194); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30874 = 6'h4 == state ? $signed(digest_47) : $signed(_GEN_30195); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30875 = 6'h4 == state ? $signed(digest_48) : $signed(_GEN_30196); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30876 = 6'h4 == state ? $signed(digest_49) : $signed(_GEN_30197); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30877 = 6'h4 == state ? $signed(digest_50) : $signed(_GEN_30198); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30878 = 6'h4 == state ? $signed(digest_51) : $signed(_GEN_30199); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30879 = 6'h4 == state ? $signed(digest_52) : $signed(_GEN_30200); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30880 = 6'h4 == state ? $signed(digest_53) : $signed(_GEN_30201); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30881 = 6'h4 == state ? $signed(digest_54) : $signed(_GEN_30202); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30882 = 6'h4 == state ? $signed(digest_55) : $signed(_GEN_30203); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30883 = 6'h4 == state ? $signed(digest_56) : $signed(_GEN_30204); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30884 = 6'h4 == state ? $signed(digest_57) : $signed(_GEN_30205); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30885 = 6'h4 == state ? $signed(digest_58) : $signed(_GEN_30206); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30886 = 6'h4 == state ? $signed(digest_59) : $signed(_GEN_30207); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30887 = 6'h4 == state ? $signed(digest_60) : $signed(_GEN_30208); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30888 = 6'h4 == state ? $signed(digest_61) : $signed(_GEN_30209); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30889 = 6'h4 == state ? $signed(digest_62) : $signed(_GEN_30210); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30890 = 6'h4 == state ? $signed(digest_63) : $signed(_GEN_30211); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30891 = 6'h4 == state ? $signed(digest_64) : $signed(_GEN_30212); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30892 = 6'h4 == state ? $signed(digest_65) : $signed(_GEN_30213); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30893 = 6'h4 == state ? $signed(digest_66) : $signed(_GEN_30214); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30894 = 6'h4 == state ? $signed(digest_67) : $signed(_GEN_30215); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30895 = 6'h4 == state ? $signed(digest_68) : $signed(_GEN_30216); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30896 = 6'h4 == state ? $signed(digest_69) : $signed(_GEN_30217); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30897 = 6'h4 == state ? $signed(digest_70) : $signed(_GEN_30218); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30898 = 6'h4 == state ? $signed(digest_71) : $signed(_GEN_30219); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30899 = 6'h4 == state ? $signed(digest_72) : $signed(_GEN_30220); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30900 = 6'h4 == state ? $signed(digest_73) : $signed(_GEN_30221); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30901 = 6'h4 == state ? $signed(digest_74) : $signed(_GEN_30222); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30902 = 6'h4 == state ? $signed(digest_75) : $signed(_GEN_30223); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30903 = 6'h4 == state ? $signed(digest_76) : $signed(_GEN_30224); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30904 = 6'h4 == state ? $signed(digest_77) : $signed(_GEN_30225); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30905 = 6'h4 == state ? $signed(digest_78) : $signed(_GEN_30226); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_30906 = 6'h4 == state ? $signed(digest_79) : $signed(_GEN_30227); // @[digest.scala 81:19 53:21]
  wire  _GEN_30908 = 6'h4 == state ? 1'h0 : _GEN_30229; // @[digest.scala 81:19 58:25]
  wire  _GEN_30991 = 6'h4 == state ? 1'h0 : _GEN_30312; // @[digest.scala 81:19 63:25]
  wire  _GEN_31074 = 6'h4 == state ? 1'h0 : _GEN_30395; // @[digest.scala 81:19 68:25]
  wire  _GEN_31157 = 6'h4 == state ? 1'h0 : _GEN_30478; // @[digest.scala 81:19 73:25]
  wire  _GEN_31240 = 6'h4 == state ? 1'h0 : _GEN_30561; // @[digest.scala 81:19 78:25]
  wire [5:0] _GEN_31241 = 6'h3 == state ? {{3'd0}, _state_T_2} : _GEN_30563; // @[digest.scala 81:19 98:19]
  wire [62:0] _GEN_31242 = 6'h3 == state ? $signed({{31{temp[31]}},temp}) : $signed(_GEN_30562); // @[digest.scala 38:19 81:19]
  wire [31:0] _GEN_31243 = 6'h3 == state ? $signed(blks_0) : $signed(_GEN_30564); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31244 = 6'h3 == state ? $signed(blks_1) : $signed(_GEN_30565); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31245 = 6'h3 == state ? $signed(blks_2) : $signed(_GEN_30566); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31246 = 6'h3 == state ? $signed(blks_3) : $signed(_GEN_30567); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31247 = 6'h3 == state ? $signed(blks_4) : $signed(_GEN_30568); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31248 = 6'h3 == state ? $signed(blks_5) : $signed(_GEN_30569); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31249 = 6'h3 == state ? $signed(blks_6) : $signed(_GEN_30570); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31250 = 6'h3 == state ? $signed(blks_7) : $signed(_GEN_30571); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31251 = 6'h3 == state ? $signed(blks_8) : $signed(_GEN_30572); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31252 = 6'h3 == state ? $signed(blks_9) : $signed(_GEN_30573); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31253 = 6'h3 == state ? $signed(blks_10) : $signed(_GEN_30574); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31254 = 6'h3 == state ? $signed(blks_11) : $signed(_GEN_30575); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31255 = 6'h3 == state ? $signed(blks_12) : $signed(_GEN_30576); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31256 = 6'h3 == state ? $signed(blks_13) : $signed(_GEN_30577); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31257 = 6'h3 == state ? $signed(blks_14) : $signed(_GEN_30578); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31258 = 6'h3 == state ? $signed(blks_15) : $signed(_GEN_30579); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31259 = 6'h3 == state ? $signed(blks_16) : $signed(_GEN_30580); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31260 = 6'h3 == state ? $signed(blks_17) : $signed(_GEN_30581); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31261 = 6'h3 == state ? $signed(blks_18) : $signed(_GEN_30582); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31262 = 6'h3 == state ? $signed(blks_19) : $signed(_GEN_30583); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31263 = 6'h3 == state ? $signed(blks_20) : $signed(_GEN_30584); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31264 = 6'h3 == state ? $signed(blks_21) : $signed(_GEN_30585); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31265 = 6'h3 == state ? $signed(blks_22) : $signed(_GEN_30586); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31266 = 6'h3 == state ? $signed(blks_23) : $signed(_GEN_30587); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31267 = 6'h3 == state ? $signed(blks_24) : $signed(_GEN_30588); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31268 = 6'h3 == state ? $signed(blks_25) : $signed(_GEN_30589); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31269 = 6'h3 == state ? $signed(blks_26) : $signed(_GEN_30590); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31270 = 6'h3 == state ? $signed(blks_27) : $signed(_GEN_30591); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31271 = 6'h3 == state ? $signed(blks_28) : $signed(_GEN_30592); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31272 = 6'h3 == state ? $signed(blks_29) : $signed(_GEN_30593); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31273 = 6'h3 == state ? $signed(blks_30) : $signed(_GEN_30594); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31274 = 6'h3 == state ? $signed(blks_31) : $signed(_GEN_30595); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31275 = 6'h3 == state ? $signed(blks_32) : $signed(_GEN_30596); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31276 = 6'h3 == state ? $signed(blks_33) : $signed(_GEN_30597); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31277 = 6'h3 == state ? $signed(blks_34) : $signed(_GEN_30598); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31278 = 6'h3 == state ? $signed(blks_35) : $signed(_GEN_30599); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31279 = 6'h3 == state ? $signed(blks_36) : $signed(_GEN_30600); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31280 = 6'h3 == state ? $signed(blks_37) : $signed(_GEN_30601); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31281 = 6'h3 == state ? $signed(blks_38) : $signed(_GEN_30602); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31282 = 6'h3 == state ? $signed(blks_39) : $signed(_GEN_30603); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31283 = 6'h3 == state ? $signed(blks_40) : $signed(_GEN_30604); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31284 = 6'h3 == state ? $signed(blks_41) : $signed(_GEN_30605); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31285 = 6'h3 == state ? $signed(blks_42) : $signed(_GEN_30606); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31286 = 6'h3 == state ? $signed(blks_43) : $signed(_GEN_30607); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31287 = 6'h3 == state ? $signed(blks_44) : $signed(_GEN_30608); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31288 = 6'h3 == state ? $signed(blks_45) : $signed(_GEN_30609); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31289 = 6'h3 == state ? $signed(blks_46) : $signed(_GEN_30610); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31290 = 6'h3 == state ? $signed(blks_47) : $signed(_GEN_30611); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31291 = 6'h3 == state ? $signed(blks_48) : $signed(_GEN_30612); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31292 = 6'h3 == state ? $signed(blks_49) : $signed(_GEN_30613); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31293 = 6'h3 == state ? $signed(blks_50) : $signed(_GEN_30614); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31294 = 6'h3 == state ? $signed(blks_51) : $signed(_GEN_30615); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31295 = 6'h3 == state ? $signed(blks_52) : $signed(_GEN_30616); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31296 = 6'h3 == state ? $signed(blks_53) : $signed(_GEN_30617); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31297 = 6'h3 == state ? $signed(blks_54) : $signed(_GEN_30618); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31298 = 6'h3 == state ? $signed(blks_55) : $signed(_GEN_30619); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31299 = 6'h3 == state ? $signed(blks_56) : $signed(_GEN_30620); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31300 = 6'h3 == state ? $signed(blks_57) : $signed(_GEN_30621); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31301 = 6'h3 == state ? $signed(blks_58) : $signed(_GEN_30622); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31302 = 6'h3 == state ? $signed(blks_59) : $signed(_GEN_30623); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31303 = 6'h3 == state ? $signed(blks_60) : $signed(_GEN_30624); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31304 = 6'h3 == state ? $signed(blks_61) : $signed(_GEN_30625); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31305 = 6'h3 == state ? $signed(blks_62) : $signed(_GEN_30626); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31306 = 6'h3 == state ? $signed(blks_63) : $signed(_GEN_30627); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31307 = 6'h3 == state ? $signed(blks_64) : $signed(_GEN_30628); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31308 = 6'h3 == state ? $signed(blks_65) : $signed(_GEN_30629); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31309 = 6'h3 == state ? $signed(blks_66) : $signed(_GEN_30630); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31310 = 6'h3 == state ? $signed(blks_67) : $signed(_GEN_30631); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31311 = 6'h3 == state ? $signed(blks_68) : $signed(_GEN_30632); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31312 = 6'h3 == state ? $signed(blks_69) : $signed(_GEN_30633); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31313 = 6'h3 == state ? $signed(blks_70) : $signed(_GEN_30634); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31314 = 6'h3 == state ? $signed(blks_71) : $signed(_GEN_30635); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31315 = 6'h3 == state ? $signed(blks_72) : $signed(_GEN_30636); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31316 = 6'h3 == state ? $signed(blks_73) : $signed(_GEN_30637); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31317 = 6'h3 == state ? $signed(blks_74) : $signed(_GEN_30638); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31318 = 6'h3 == state ? $signed(blks_75) : $signed(_GEN_30639); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31319 = 6'h3 == state ? $signed(blks_76) : $signed(_GEN_30640); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31320 = 6'h3 == state ? $signed(blks_77) : $signed(_GEN_30641); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31321 = 6'h3 == state ? $signed(blks_78) : $signed(_GEN_30642); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31322 = 6'h3 == state ? $signed(blks_79) : $signed(_GEN_30643); // @[digest.scala 39:19 81:19]
  wire [31:0] _GEN_31323 = 6'h3 == state ? $signed(i) : $signed(_GEN_30644); // @[digest.scala 23:16 81:19]
  wire [31:0] _GEN_31324 = 6'h3 == state ? $signed(a) : $signed(_GEN_30645); // @[digest.scala 24:16 81:19]
  wire [31:0] _GEN_31325 = 6'h3 == state ? $signed(b) : $signed(_GEN_30646); // @[digest.scala 25:16 81:19]
  wire [31:0] _GEN_31326 = 6'h3 == state ? $signed(c) : $signed(_GEN_30647); // @[digest.scala 26:16 81:19]
  wire [31:0] _GEN_31327 = 6'h3 == state ? $signed(d) : $signed(_GEN_30648); // @[digest.scala 27:16 81:19]
  wire [31:0] _GEN_31328 = 6'h3 == state ? $signed(e) : $signed(_GEN_30649); // @[digest.scala 28:16 81:19]
  wire [31:0] _GEN_31329 = 6'h3 == state ? $signed(olda) : $signed(_GEN_30650); // @[digest.scala 29:19 81:19]
  wire [31:0] _GEN_31330 = 6'h3 == state ? $signed(oldb) : $signed(_GEN_30651); // @[digest.scala 30:19 81:19]
  wire [31:0] _GEN_31331 = 6'h3 == state ? $signed(oldc) : $signed(_GEN_30652); // @[digest.scala 31:19 81:19]
  wire [31:0] _GEN_31332 = 6'h3 == state ? $signed(oldd) : $signed(_GEN_30653); // @[digest.scala 32:19 81:19]
  wire [31:0] _GEN_31333 = 6'h3 == state ? $signed(olde) : $signed(_GEN_30654); // @[digest.scala 33:19 81:19]
  wire [31:0] _GEN_31334 = 6'h3 == state ? $signed(j) : $signed(_GEN_30655); // @[digest.scala 34:16 81:19]
  wire [31:0] _GEN_31335 = 6'h3 == state ? $signed(w_0) : $signed(_GEN_30656); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31336 = 6'h3 == state ? $signed(w_1) : $signed(_GEN_30657); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31337 = 6'h3 == state ? $signed(w_2) : $signed(_GEN_30658); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31338 = 6'h3 == state ? $signed(w_3) : $signed(_GEN_30659); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31339 = 6'h3 == state ? $signed(w_4) : $signed(_GEN_30660); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31340 = 6'h3 == state ? $signed(w_5) : $signed(_GEN_30661); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31341 = 6'h3 == state ? $signed(w_6) : $signed(_GEN_30662); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31342 = 6'h3 == state ? $signed(w_7) : $signed(_GEN_30663); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31343 = 6'h3 == state ? $signed(w_8) : $signed(_GEN_30664); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31344 = 6'h3 == state ? $signed(w_9) : $signed(_GEN_30665); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31345 = 6'h3 == state ? $signed(w_10) : $signed(_GEN_30666); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31346 = 6'h3 == state ? $signed(w_11) : $signed(_GEN_30667); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31347 = 6'h3 == state ? $signed(w_12) : $signed(_GEN_30668); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31348 = 6'h3 == state ? $signed(w_13) : $signed(_GEN_30669); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31349 = 6'h3 == state ? $signed(w_14) : $signed(_GEN_30670); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31350 = 6'h3 == state ? $signed(w_15) : $signed(_GEN_30671); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31351 = 6'h3 == state ? $signed(w_16) : $signed(_GEN_30672); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31352 = 6'h3 == state ? $signed(w_17) : $signed(_GEN_30673); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31353 = 6'h3 == state ? $signed(w_18) : $signed(_GEN_30674); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31354 = 6'h3 == state ? $signed(w_19) : $signed(_GEN_30675); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31355 = 6'h3 == state ? $signed(w_20) : $signed(_GEN_30676); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31356 = 6'h3 == state ? $signed(w_21) : $signed(_GEN_30677); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31357 = 6'h3 == state ? $signed(w_22) : $signed(_GEN_30678); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31358 = 6'h3 == state ? $signed(w_23) : $signed(_GEN_30679); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31359 = 6'h3 == state ? $signed(w_24) : $signed(_GEN_30680); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31360 = 6'h3 == state ? $signed(w_25) : $signed(_GEN_30681); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31361 = 6'h3 == state ? $signed(w_26) : $signed(_GEN_30682); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31362 = 6'h3 == state ? $signed(w_27) : $signed(_GEN_30683); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31363 = 6'h3 == state ? $signed(w_28) : $signed(_GEN_30684); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31364 = 6'h3 == state ? $signed(w_29) : $signed(_GEN_30685); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31365 = 6'h3 == state ? $signed(w_30) : $signed(_GEN_30686); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31366 = 6'h3 == state ? $signed(w_31) : $signed(_GEN_30687); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31367 = 6'h3 == state ? $signed(w_32) : $signed(_GEN_30688); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31368 = 6'h3 == state ? $signed(w_33) : $signed(_GEN_30689); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31369 = 6'h3 == state ? $signed(w_34) : $signed(_GEN_30690); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31370 = 6'h3 == state ? $signed(w_35) : $signed(_GEN_30691); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31371 = 6'h3 == state ? $signed(w_36) : $signed(_GEN_30692); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31372 = 6'h3 == state ? $signed(w_37) : $signed(_GEN_30693); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31373 = 6'h3 == state ? $signed(w_38) : $signed(_GEN_30694); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31374 = 6'h3 == state ? $signed(w_39) : $signed(_GEN_30695); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31375 = 6'h3 == state ? $signed(w_40) : $signed(_GEN_30696); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31376 = 6'h3 == state ? $signed(w_41) : $signed(_GEN_30697); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31377 = 6'h3 == state ? $signed(w_42) : $signed(_GEN_30698); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31378 = 6'h3 == state ? $signed(w_43) : $signed(_GEN_30699); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31379 = 6'h3 == state ? $signed(w_44) : $signed(_GEN_30700); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31380 = 6'h3 == state ? $signed(w_45) : $signed(_GEN_30701); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31381 = 6'h3 == state ? $signed(w_46) : $signed(_GEN_30702); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31382 = 6'h3 == state ? $signed(w_47) : $signed(_GEN_30703); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31383 = 6'h3 == state ? $signed(w_48) : $signed(_GEN_30704); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31384 = 6'h3 == state ? $signed(w_49) : $signed(_GEN_30705); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31385 = 6'h3 == state ? $signed(w_50) : $signed(_GEN_30706); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31386 = 6'h3 == state ? $signed(w_51) : $signed(_GEN_30707); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31387 = 6'h3 == state ? $signed(w_52) : $signed(_GEN_30708); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31388 = 6'h3 == state ? $signed(w_53) : $signed(_GEN_30709); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31389 = 6'h3 == state ? $signed(w_54) : $signed(_GEN_30710); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31390 = 6'h3 == state ? $signed(w_55) : $signed(_GEN_30711); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31391 = 6'h3 == state ? $signed(w_56) : $signed(_GEN_30712); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31392 = 6'h3 == state ? $signed(w_57) : $signed(_GEN_30713); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31393 = 6'h3 == state ? $signed(w_58) : $signed(_GEN_30714); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31394 = 6'h3 == state ? $signed(w_59) : $signed(_GEN_30715); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31395 = 6'h3 == state ? $signed(w_60) : $signed(_GEN_30716); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31396 = 6'h3 == state ? $signed(w_61) : $signed(_GEN_30717); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31397 = 6'h3 == state ? $signed(w_62) : $signed(_GEN_30718); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31398 = 6'h3 == state ? $signed(w_63) : $signed(_GEN_30719); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31399 = 6'h3 == state ? $signed(w_64) : $signed(_GEN_30720); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31400 = 6'h3 == state ? $signed(w_65) : $signed(_GEN_30721); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31401 = 6'h3 == state ? $signed(w_66) : $signed(_GEN_30722); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31402 = 6'h3 == state ? $signed(w_67) : $signed(_GEN_30723); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31403 = 6'h3 == state ? $signed(w_68) : $signed(_GEN_30724); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31404 = 6'h3 == state ? $signed(w_69) : $signed(_GEN_30725); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31405 = 6'h3 == state ? $signed(w_70) : $signed(_GEN_30726); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31406 = 6'h3 == state ? $signed(w_71) : $signed(_GEN_30727); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31407 = 6'h3 == state ? $signed(w_72) : $signed(_GEN_30728); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31408 = 6'h3 == state ? $signed(w_73) : $signed(_GEN_30729); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31409 = 6'h3 == state ? $signed(w_74) : $signed(_GEN_30730); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31410 = 6'h3 == state ? $signed(w_75) : $signed(_GEN_30731); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31411 = 6'h3 == state ? $signed(w_76) : $signed(_GEN_30732); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31412 = 6'h3 == state ? $signed(w_77) : $signed(_GEN_30733); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31413 = 6'h3 == state ? $signed(w_78) : $signed(_GEN_30734); // @[digest.scala 40:16 81:19]
  wire [31:0] _GEN_31414 = 6'h3 == state ? $signed(w_79) : $signed(_GEN_30735); // @[digest.scala 40:16 81:19]
  wire  _GEN_31415 = 6'h3 == state ? 1'h0 : _GEN_30736; // @[digest.scala 81:19 44:24]
  wire [31:0] _GEN_31418 = 6'h3 == state ? $signed(t) : $signed(_GEN_30739); // @[digest.scala 35:16 81:19]
  wire  _GEN_31419 = 6'h3 == state ? 1'h0 : _GEN_30740; // @[digest.scala 81:19 48:24]
  wire  _GEN_31422 = 6'h3 == state ? 1'h0 : _GEN_30743; // @[digest.scala 81:19 52:24]
  wire [31:0] _GEN_31506 = 6'h3 == state ? $signed(digest_0) : $signed(_GEN_30827); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31507 = 6'h3 == state ? $signed(digest_1) : $signed(_GEN_30828); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31508 = 6'h3 == state ? $signed(digest_2) : $signed(_GEN_30829); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31509 = 6'h3 == state ? $signed(digest_3) : $signed(_GEN_30830); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31510 = 6'h3 == state ? $signed(digest_4) : $signed(_GEN_30831); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31511 = 6'h3 == state ? $signed(digest_5) : $signed(_GEN_30832); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31512 = 6'h3 == state ? $signed(digest_6) : $signed(_GEN_30833); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31513 = 6'h3 == state ? $signed(digest_7) : $signed(_GEN_30834); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31514 = 6'h3 == state ? $signed(digest_8) : $signed(_GEN_30835); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31515 = 6'h3 == state ? $signed(digest_9) : $signed(_GEN_30836); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31516 = 6'h3 == state ? $signed(digest_10) : $signed(_GEN_30837); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31517 = 6'h3 == state ? $signed(digest_11) : $signed(_GEN_30838); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31518 = 6'h3 == state ? $signed(digest_12) : $signed(_GEN_30839); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31519 = 6'h3 == state ? $signed(digest_13) : $signed(_GEN_30840); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31520 = 6'h3 == state ? $signed(digest_14) : $signed(_GEN_30841); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31521 = 6'h3 == state ? $signed(digest_15) : $signed(_GEN_30842); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31522 = 6'h3 == state ? $signed(digest_16) : $signed(_GEN_30843); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31523 = 6'h3 == state ? $signed(digest_17) : $signed(_GEN_30844); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31524 = 6'h3 == state ? $signed(digest_18) : $signed(_GEN_30845); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31525 = 6'h3 == state ? $signed(digest_19) : $signed(_GEN_30846); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31526 = 6'h3 == state ? $signed(digest_20) : $signed(_GEN_30847); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31527 = 6'h3 == state ? $signed(digest_21) : $signed(_GEN_30848); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31528 = 6'h3 == state ? $signed(digest_22) : $signed(_GEN_30849); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31529 = 6'h3 == state ? $signed(digest_23) : $signed(_GEN_30850); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31530 = 6'h3 == state ? $signed(digest_24) : $signed(_GEN_30851); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31531 = 6'h3 == state ? $signed(digest_25) : $signed(_GEN_30852); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31532 = 6'h3 == state ? $signed(digest_26) : $signed(_GEN_30853); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31533 = 6'h3 == state ? $signed(digest_27) : $signed(_GEN_30854); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31534 = 6'h3 == state ? $signed(digest_28) : $signed(_GEN_30855); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31535 = 6'h3 == state ? $signed(digest_29) : $signed(_GEN_30856); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31536 = 6'h3 == state ? $signed(digest_30) : $signed(_GEN_30857); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31537 = 6'h3 == state ? $signed(digest_31) : $signed(_GEN_30858); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31538 = 6'h3 == state ? $signed(digest_32) : $signed(_GEN_30859); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31539 = 6'h3 == state ? $signed(digest_33) : $signed(_GEN_30860); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31540 = 6'h3 == state ? $signed(digest_34) : $signed(_GEN_30861); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31541 = 6'h3 == state ? $signed(digest_35) : $signed(_GEN_30862); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31542 = 6'h3 == state ? $signed(digest_36) : $signed(_GEN_30863); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31543 = 6'h3 == state ? $signed(digest_37) : $signed(_GEN_30864); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31544 = 6'h3 == state ? $signed(digest_38) : $signed(_GEN_30865); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31545 = 6'h3 == state ? $signed(digest_39) : $signed(_GEN_30866); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31546 = 6'h3 == state ? $signed(digest_40) : $signed(_GEN_30867); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31547 = 6'h3 == state ? $signed(digest_41) : $signed(_GEN_30868); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31548 = 6'h3 == state ? $signed(digest_42) : $signed(_GEN_30869); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31549 = 6'h3 == state ? $signed(digest_43) : $signed(_GEN_30870); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31550 = 6'h3 == state ? $signed(digest_44) : $signed(_GEN_30871); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31551 = 6'h3 == state ? $signed(digest_45) : $signed(_GEN_30872); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31552 = 6'h3 == state ? $signed(digest_46) : $signed(_GEN_30873); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31553 = 6'h3 == state ? $signed(digest_47) : $signed(_GEN_30874); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31554 = 6'h3 == state ? $signed(digest_48) : $signed(_GEN_30875); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31555 = 6'h3 == state ? $signed(digest_49) : $signed(_GEN_30876); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31556 = 6'h3 == state ? $signed(digest_50) : $signed(_GEN_30877); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31557 = 6'h3 == state ? $signed(digest_51) : $signed(_GEN_30878); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31558 = 6'h3 == state ? $signed(digest_52) : $signed(_GEN_30879); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31559 = 6'h3 == state ? $signed(digest_53) : $signed(_GEN_30880); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31560 = 6'h3 == state ? $signed(digest_54) : $signed(_GEN_30881); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31561 = 6'h3 == state ? $signed(digest_55) : $signed(_GEN_30882); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31562 = 6'h3 == state ? $signed(digest_56) : $signed(_GEN_30883); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31563 = 6'h3 == state ? $signed(digest_57) : $signed(_GEN_30884); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31564 = 6'h3 == state ? $signed(digest_58) : $signed(_GEN_30885); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31565 = 6'h3 == state ? $signed(digest_59) : $signed(_GEN_30886); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31566 = 6'h3 == state ? $signed(digest_60) : $signed(_GEN_30887); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31567 = 6'h3 == state ? $signed(digest_61) : $signed(_GEN_30888); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31568 = 6'h3 == state ? $signed(digest_62) : $signed(_GEN_30889); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31569 = 6'h3 == state ? $signed(digest_63) : $signed(_GEN_30890); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31570 = 6'h3 == state ? $signed(digest_64) : $signed(_GEN_30891); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31571 = 6'h3 == state ? $signed(digest_65) : $signed(_GEN_30892); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31572 = 6'h3 == state ? $signed(digest_66) : $signed(_GEN_30893); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31573 = 6'h3 == state ? $signed(digest_67) : $signed(_GEN_30894); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31574 = 6'h3 == state ? $signed(digest_68) : $signed(_GEN_30895); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31575 = 6'h3 == state ? $signed(digest_69) : $signed(_GEN_30896); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31576 = 6'h3 == state ? $signed(digest_70) : $signed(_GEN_30897); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31577 = 6'h3 == state ? $signed(digest_71) : $signed(_GEN_30898); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31578 = 6'h3 == state ? $signed(digest_72) : $signed(_GEN_30899); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31579 = 6'h3 == state ? $signed(digest_73) : $signed(_GEN_30900); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31580 = 6'h3 == state ? $signed(digest_74) : $signed(_GEN_30901); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31581 = 6'h3 == state ? $signed(digest_75) : $signed(_GEN_30902); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31582 = 6'h3 == state ? $signed(digest_76) : $signed(_GEN_30903); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31583 = 6'h3 == state ? $signed(digest_77) : $signed(_GEN_30904); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31584 = 6'h3 == state ? $signed(digest_78) : $signed(_GEN_30905); // @[digest.scala 81:19 53:21]
  wire [31:0] _GEN_31585 = 6'h3 == state ? $signed(digest_79) : $signed(_GEN_30906); // @[digest.scala 81:19 53:21]
  wire  _GEN_31587 = 6'h3 == state ? 1'h0 : _GEN_30908; // @[digest.scala 81:19 58:25]
  wire  _GEN_31670 = 6'h3 == state ? 1'h0 : _GEN_30991; // @[digest.scala 81:19 63:25]
  wire  _GEN_31753 = 6'h3 == state ? 1'h0 : _GEN_31074; // @[digest.scala 81:19 68:25]
  wire  _GEN_31836 = 6'h3 == state ? 1'h0 : _GEN_31157; // @[digest.scala 81:19 73:25]
  wire  _GEN_31919 = 6'h3 == state ? 1'h0 : _GEN_31240; // @[digest.scala 81:19 78:25]
  wire [5:0] _GEN_31921 = 6'h2 == state ? 6'h3 : _GEN_31241; // @[digest.scala 81:19 95:19]
  wire [62:0] _GEN_31922 = 6'h2 == state ? $signed({{31{temp[31]}},temp}) : $signed(_GEN_31242); // @[digest.scala 38:19 81:19]
  wire  _GEN_32094 = 6'h2 == state ? 1'h0 : _GEN_31415; // @[digest.scala 81:19 44:24]
  wire  _GEN_32098 = 6'h2 == state ? 1'h0 : _GEN_31419; // @[digest.scala 81:19 48:24]
  wire  _GEN_32101 = 6'h2 == state ? 1'h0 : _GEN_31422; // @[digest.scala 81:19 52:24]
  wire  _GEN_32266 = 6'h2 == state ? 1'h0 : _GEN_31587; // @[digest.scala 81:19 58:25]
  wire  _GEN_32349 = 6'h2 == state ? 1'h0 : _GEN_31670; // @[digest.scala 81:19 63:25]
  wire  _GEN_32432 = 6'h2 == state ? 1'h0 : _GEN_31753; // @[digest.scala 81:19 68:25]
  wire  _GEN_32515 = 6'h2 == state ? 1'h0 : _GEN_31836; // @[digest.scala 81:19 73:25]
  wire  _GEN_32598 = 6'h2 == state ? 1'h0 : _GEN_31919; // @[digest.scala 81:19 78:25]
  wire [63:0] _GEN_32599 = 6'h1 == state ? $signed(_blksLength_T_9) : $signed({{32{blksLength[31]}},blksLength}); // @[digest.scala 81:19 90:24 37:25]
  wire [62:0] _GEN_32602 = 6'h1 == state ? $signed({{31{temp[31]}},temp}) : $signed(_GEN_31922); // @[digest.scala 38:19 81:19]
  wire  _GEN_32774 = 6'h1 == state ? 1'h0 : _GEN_32094; // @[digest.scala 81:19 44:24]
  wire  _GEN_32778 = 6'h1 == state ? 1'h0 : _GEN_32098; // @[digest.scala 81:19 48:24]
  wire  _GEN_32781 = 6'h1 == state ? 1'h0 : _GEN_32101; // @[digest.scala 81:19 52:24]
  wire  _GEN_32946 = 6'h1 == state ? 1'h0 : _GEN_32266; // @[digest.scala 81:19 58:25]
  wire  _GEN_33029 = 6'h1 == state ? 1'h0 : _GEN_32349; // @[digest.scala 81:19 63:25]
  wire  _GEN_33112 = 6'h1 == state ? 1'h0 : _GEN_32432; // @[digest.scala 81:19 68:25]
  wire  _GEN_33195 = 6'h1 == state ? 1'h0 : _GEN_32515; // @[digest.scala 81:19 73:25]
  wire  _GEN_33278 = 6'h1 == state ? 1'h0 : _GEN_32598; // @[digest.scala 81:19 78:25]
  wire [63:0] _GEN_33281 = 6'h0 == state ? $signed({{32{blksLength[31]}},blksLength}) : $signed(_GEN_32599); // @[digest.scala 81:19 37:25]
  wire [62:0] _GEN_33283 = 6'h0 == state ? $signed({{31{temp[31]}},temp}) : $signed(_GEN_32602); // @[digest.scala 38:19 81:19]
  wire  _GEN_33455 = 6'h0 == state ? 1'h0 : _GEN_32774; // @[digest.scala 81:19 44:24]
  wire  _GEN_33459 = 6'h0 == state ? 1'h0 : _GEN_32778; // @[digest.scala 81:19 48:24]
  wire  _GEN_33462 = 6'h0 == state ? 1'h0 : _GEN_32781; // @[digest.scala 81:19 52:24]
  wire  _GEN_33627 = 6'h0 == state ? 1'h0 : _GEN_32946; // @[digest.scala 81:19 58:25]
  wire  _GEN_33710 = 6'h0 == state ? 1'h0 : _GEN_33029; // @[digest.scala 81:19 63:25]
  wire  _GEN_33793 = 6'h0 == state ? 1'h0 : _GEN_33112; // @[digest.scala 81:19 68:25]
  wire  _GEN_33876 = 6'h0 == state ? 1'h0 : _GEN_33195; // @[digest.scala 81:19 73:25]
  wire  _GEN_33959 = 6'h0 == state ? 1'h0 : _GEN_33278; // @[digest.scala 81:19 78:25]
  wire [63:0] _GEN_33962 = 6'h3f == state ? $signed({{32{blksLength[31]}},blksLength}) : $signed(_GEN_33281); // @[digest.scala 81:19 37:25]
  wire [62:0] _GEN_33964 = 6'h3f == state ? $signed({{31{temp[31]}},temp}) : $signed(_GEN_33283); // @[digest.scala 38:19 81:19]
  rol __m_rol_0 ( // @[digest.scala 41:27]
    .clock(__m_rol_0_clock),
    .reset(__m_rol_0_reset),
    .io_num(__m_rol_0_io_num),
    .io_cnt(__m_rol_0_io_cnt),
    .io_valid(__m_rol_0_io_valid),
    .io_ready(__m_rol_0_io_ready),
    .io_out_rol(__m_rol_0_io_out_rol)
  );
  rol __m_rol_1 ( // @[digest.scala 45:27]
    .clock(__m_rol_1_clock),
    .reset(__m_rol_1_reset),
    .io_num(__m_rol_1_io_num),
    .io_cnt(__m_rol_1_io_cnt),
    .io_valid(__m_rol_1_io_valid),
    .io_ready(__m_rol_1_io_ready),
    .io_out_rol(__m_rol_1_io_out_rol)
  );
  rol __m_rol_2 ( // @[digest.scala 49:27]
    .clock(__m_rol_2_clock),
    .reset(__m_rol_2_reset),
    .io_num(__m_rol_2_io_num),
    .io_cnt(__m_rol_2_io_cnt),
    .io_valid(__m_rol_2_io_valid),
    .io_ready(__m_rol_2_io_ready),
    .io_out_rol(__m_rol_2_io_out_rol)
  );
  fill __m_fill_0 ( // @[digest.scala 54:28]
    .clock(__m_fill_0_clock),
    .reset(__m_fill_0_reset),
    .io_value(__m_fill_0_io_value),
    .io_arr_0(__m_fill_0_io_arr_0),
    .io_arr_1(__m_fill_0_io_arr_1),
    .io_arr_2(__m_fill_0_io_arr_2),
    .io_arr_3(__m_fill_0_io_arr_3),
    .io_arr_4(__m_fill_0_io_arr_4),
    .io_arr_5(__m_fill_0_io_arr_5),
    .io_arr_6(__m_fill_0_io_arr_6),
    .io_arr_7(__m_fill_0_io_arr_7),
    .io_arr_8(__m_fill_0_io_arr_8),
    .io_arr_9(__m_fill_0_io_arr_9),
    .io_arr_10(__m_fill_0_io_arr_10),
    .io_arr_11(__m_fill_0_io_arr_11),
    .io_arr_12(__m_fill_0_io_arr_12),
    .io_arr_13(__m_fill_0_io_arr_13),
    .io_arr_14(__m_fill_0_io_arr_14),
    .io_arr_15(__m_fill_0_io_arr_15),
    .io_arr_16(__m_fill_0_io_arr_16),
    .io_arr_17(__m_fill_0_io_arr_17),
    .io_arr_18(__m_fill_0_io_arr_18),
    .io_arr_19(__m_fill_0_io_arr_19),
    .io_arr_20(__m_fill_0_io_arr_20),
    .io_arr_21(__m_fill_0_io_arr_21),
    .io_arr_22(__m_fill_0_io_arr_22),
    .io_arr_23(__m_fill_0_io_arr_23),
    .io_arr_24(__m_fill_0_io_arr_24),
    .io_arr_25(__m_fill_0_io_arr_25),
    .io_arr_26(__m_fill_0_io_arr_26),
    .io_arr_27(__m_fill_0_io_arr_27),
    .io_arr_28(__m_fill_0_io_arr_28),
    .io_arr_29(__m_fill_0_io_arr_29),
    .io_arr_30(__m_fill_0_io_arr_30),
    .io_arr_31(__m_fill_0_io_arr_31),
    .io_arr_32(__m_fill_0_io_arr_32),
    .io_arr_33(__m_fill_0_io_arr_33),
    .io_arr_34(__m_fill_0_io_arr_34),
    .io_arr_35(__m_fill_0_io_arr_35),
    .io_arr_36(__m_fill_0_io_arr_36),
    .io_arr_37(__m_fill_0_io_arr_37),
    .io_arr_38(__m_fill_0_io_arr_38),
    .io_arr_39(__m_fill_0_io_arr_39),
    .io_arr_40(__m_fill_0_io_arr_40),
    .io_arr_41(__m_fill_0_io_arr_41),
    .io_arr_42(__m_fill_0_io_arr_42),
    .io_arr_43(__m_fill_0_io_arr_43),
    .io_arr_44(__m_fill_0_io_arr_44),
    .io_arr_45(__m_fill_0_io_arr_45),
    .io_arr_46(__m_fill_0_io_arr_46),
    .io_arr_47(__m_fill_0_io_arr_47),
    .io_arr_48(__m_fill_0_io_arr_48),
    .io_arr_49(__m_fill_0_io_arr_49),
    .io_arr_50(__m_fill_0_io_arr_50),
    .io_arr_51(__m_fill_0_io_arr_51),
    .io_arr_52(__m_fill_0_io_arr_52),
    .io_arr_53(__m_fill_0_io_arr_53),
    .io_arr_54(__m_fill_0_io_arr_54),
    .io_arr_55(__m_fill_0_io_arr_55),
    .io_arr_56(__m_fill_0_io_arr_56),
    .io_arr_57(__m_fill_0_io_arr_57),
    .io_arr_58(__m_fill_0_io_arr_58),
    .io_arr_59(__m_fill_0_io_arr_59),
    .io_arr_60(__m_fill_0_io_arr_60),
    .io_arr_61(__m_fill_0_io_arr_61),
    .io_arr_62(__m_fill_0_io_arr_62),
    .io_arr_63(__m_fill_0_io_arr_63),
    .io_arr_64(__m_fill_0_io_arr_64),
    .io_arr_65(__m_fill_0_io_arr_65),
    .io_arr_66(__m_fill_0_io_arr_66),
    .io_arr_67(__m_fill_0_io_arr_67),
    .io_arr_68(__m_fill_0_io_arr_68),
    .io_arr_69(__m_fill_0_io_arr_69),
    .io_arr_70(__m_fill_0_io_arr_70),
    .io_arr_71(__m_fill_0_io_arr_71),
    .io_arr_72(__m_fill_0_io_arr_72),
    .io_arr_73(__m_fill_0_io_arr_73),
    .io_arr_74(__m_fill_0_io_arr_74),
    .io_arr_75(__m_fill_0_io_arr_75),
    .io_arr_76(__m_fill_0_io_arr_76),
    .io_arr_77(__m_fill_0_io_arr_77),
    .io_arr_78(__m_fill_0_io_arr_78),
    .io_arr_79(__m_fill_0_io_arr_79),
    .io_off(__m_fill_0_io_off),
    .io_valid(__m_fill_0_io_valid),
    .io_arr_out_0(__m_fill_0_io_arr_out_0),
    .io_arr_out_1(__m_fill_0_io_arr_out_1),
    .io_arr_out_2(__m_fill_0_io_arr_out_2),
    .io_arr_out_3(__m_fill_0_io_arr_out_3),
    .io_arr_out_4(__m_fill_0_io_arr_out_4),
    .io_arr_out_5(__m_fill_0_io_arr_out_5),
    .io_arr_out_6(__m_fill_0_io_arr_out_6),
    .io_arr_out_7(__m_fill_0_io_arr_out_7),
    .io_arr_out_8(__m_fill_0_io_arr_out_8),
    .io_arr_out_9(__m_fill_0_io_arr_out_9),
    .io_arr_out_10(__m_fill_0_io_arr_out_10),
    .io_arr_out_11(__m_fill_0_io_arr_out_11),
    .io_arr_out_12(__m_fill_0_io_arr_out_12),
    .io_arr_out_13(__m_fill_0_io_arr_out_13),
    .io_arr_out_14(__m_fill_0_io_arr_out_14),
    .io_arr_out_15(__m_fill_0_io_arr_out_15),
    .io_arr_out_16(__m_fill_0_io_arr_out_16),
    .io_arr_out_17(__m_fill_0_io_arr_out_17),
    .io_arr_out_18(__m_fill_0_io_arr_out_18),
    .io_arr_out_19(__m_fill_0_io_arr_out_19),
    .io_arr_out_20(__m_fill_0_io_arr_out_20),
    .io_arr_out_21(__m_fill_0_io_arr_out_21),
    .io_arr_out_22(__m_fill_0_io_arr_out_22),
    .io_arr_out_23(__m_fill_0_io_arr_out_23),
    .io_arr_out_24(__m_fill_0_io_arr_out_24),
    .io_arr_out_25(__m_fill_0_io_arr_out_25),
    .io_arr_out_26(__m_fill_0_io_arr_out_26),
    .io_arr_out_27(__m_fill_0_io_arr_out_27),
    .io_arr_out_28(__m_fill_0_io_arr_out_28),
    .io_arr_out_29(__m_fill_0_io_arr_out_29),
    .io_arr_out_30(__m_fill_0_io_arr_out_30),
    .io_arr_out_31(__m_fill_0_io_arr_out_31),
    .io_arr_out_32(__m_fill_0_io_arr_out_32),
    .io_arr_out_33(__m_fill_0_io_arr_out_33),
    .io_arr_out_34(__m_fill_0_io_arr_out_34),
    .io_arr_out_35(__m_fill_0_io_arr_out_35),
    .io_arr_out_36(__m_fill_0_io_arr_out_36),
    .io_arr_out_37(__m_fill_0_io_arr_out_37),
    .io_arr_out_38(__m_fill_0_io_arr_out_38),
    .io_arr_out_39(__m_fill_0_io_arr_out_39),
    .io_arr_out_40(__m_fill_0_io_arr_out_40),
    .io_arr_out_41(__m_fill_0_io_arr_out_41),
    .io_arr_out_42(__m_fill_0_io_arr_out_42),
    .io_arr_out_43(__m_fill_0_io_arr_out_43),
    .io_arr_out_44(__m_fill_0_io_arr_out_44),
    .io_arr_out_45(__m_fill_0_io_arr_out_45),
    .io_arr_out_46(__m_fill_0_io_arr_out_46),
    .io_arr_out_47(__m_fill_0_io_arr_out_47),
    .io_arr_out_48(__m_fill_0_io_arr_out_48),
    .io_arr_out_49(__m_fill_0_io_arr_out_49),
    .io_arr_out_50(__m_fill_0_io_arr_out_50),
    .io_arr_out_51(__m_fill_0_io_arr_out_51),
    .io_arr_out_52(__m_fill_0_io_arr_out_52),
    .io_arr_out_53(__m_fill_0_io_arr_out_53),
    .io_arr_out_54(__m_fill_0_io_arr_out_54),
    .io_arr_out_55(__m_fill_0_io_arr_out_55),
    .io_arr_out_56(__m_fill_0_io_arr_out_56),
    .io_arr_out_57(__m_fill_0_io_arr_out_57),
    .io_arr_out_58(__m_fill_0_io_arr_out_58),
    .io_arr_out_59(__m_fill_0_io_arr_out_59),
    .io_arr_out_60(__m_fill_0_io_arr_out_60),
    .io_arr_out_61(__m_fill_0_io_arr_out_61),
    .io_arr_out_62(__m_fill_0_io_arr_out_62),
    .io_arr_out_63(__m_fill_0_io_arr_out_63),
    .io_arr_out_64(__m_fill_0_io_arr_out_64),
    .io_arr_out_65(__m_fill_0_io_arr_out_65),
    .io_arr_out_66(__m_fill_0_io_arr_out_66),
    .io_arr_out_67(__m_fill_0_io_arr_out_67),
    .io_arr_out_68(__m_fill_0_io_arr_out_68),
    .io_arr_out_69(__m_fill_0_io_arr_out_69),
    .io_arr_out_70(__m_fill_0_io_arr_out_70),
    .io_arr_out_71(__m_fill_0_io_arr_out_71),
    .io_arr_out_72(__m_fill_0_io_arr_out_72),
    .io_arr_out_73(__m_fill_0_io_arr_out_73),
    .io_arr_out_74(__m_fill_0_io_arr_out_74),
    .io_arr_out_75(__m_fill_0_io_arr_out_75),
    .io_arr_out_76(__m_fill_0_io_arr_out_76),
    .io_arr_out_77(__m_fill_0_io_arr_out_77),
    .io_arr_out_78(__m_fill_0_io_arr_out_78),
    .io_arr_out_79(__m_fill_0_io_arr_out_79),
    .io_ready(__m_fill_0_io_ready)
  );
  fill __m_fill_1 ( // @[digest.scala 59:28]
    .clock(__m_fill_1_clock),
    .reset(__m_fill_1_reset),
    .io_value(__m_fill_1_io_value),
    .io_arr_0(__m_fill_1_io_arr_0),
    .io_arr_1(__m_fill_1_io_arr_1),
    .io_arr_2(__m_fill_1_io_arr_2),
    .io_arr_3(__m_fill_1_io_arr_3),
    .io_arr_4(__m_fill_1_io_arr_4),
    .io_arr_5(__m_fill_1_io_arr_5),
    .io_arr_6(__m_fill_1_io_arr_6),
    .io_arr_7(__m_fill_1_io_arr_7),
    .io_arr_8(__m_fill_1_io_arr_8),
    .io_arr_9(__m_fill_1_io_arr_9),
    .io_arr_10(__m_fill_1_io_arr_10),
    .io_arr_11(__m_fill_1_io_arr_11),
    .io_arr_12(__m_fill_1_io_arr_12),
    .io_arr_13(__m_fill_1_io_arr_13),
    .io_arr_14(__m_fill_1_io_arr_14),
    .io_arr_15(__m_fill_1_io_arr_15),
    .io_arr_16(__m_fill_1_io_arr_16),
    .io_arr_17(__m_fill_1_io_arr_17),
    .io_arr_18(__m_fill_1_io_arr_18),
    .io_arr_19(__m_fill_1_io_arr_19),
    .io_arr_20(__m_fill_1_io_arr_20),
    .io_arr_21(__m_fill_1_io_arr_21),
    .io_arr_22(__m_fill_1_io_arr_22),
    .io_arr_23(__m_fill_1_io_arr_23),
    .io_arr_24(__m_fill_1_io_arr_24),
    .io_arr_25(__m_fill_1_io_arr_25),
    .io_arr_26(__m_fill_1_io_arr_26),
    .io_arr_27(__m_fill_1_io_arr_27),
    .io_arr_28(__m_fill_1_io_arr_28),
    .io_arr_29(__m_fill_1_io_arr_29),
    .io_arr_30(__m_fill_1_io_arr_30),
    .io_arr_31(__m_fill_1_io_arr_31),
    .io_arr_32(__m_fill_1_io_arr_32),
    .io_arr_33(__m_fill_1_io_arr_33),
    .io_arr_34(__m_fill_1_io_arr_34),
    .io_arr_35(__m_fill_1_io_arr_35),
    .io_arr_36(__m_fill_1_io_arr_36),
    .io_arr_37(__m_fill_1_io_arr_37),
    .io_arr_38(__m_fill_1_io_arr_38),
    .io_arr_39(__m_fill_1_io_arr_39),
    .io_arr_40(__m_fill_1_io_arr_40),
    .io_arr_41(__m_fill_1_io_arr_41),
    .io_arr_42(__m_fill_1_io_arr_42),
    .io_arr_43(__m_fill_1_io_arr_43),
    .io_arr_44(__m_fill_1_io_arr_44),
    .io_arr_45(__m_fill_1_io_arr_45),
    .io_arr_46(__m_fill_1_io_arr_46),
    .io_arr_47(__m_fill_1_io_arr_47),
    .io_arr_48(__m_fill_1_io_arr_48),
    .io_arr_49(__m_fill_1_io_arr_49),
    .io_arr_50(__m_fill_1_io_arr_50),
    .io_arr_51(__m_fill_1_io_arr_51),
    .io_arr_52(__m_fill_1_io_arr_52),
    .io_arr_53(__m_fill_1_io_arr_53),
    .io_arr_54(__m_fill_1_io_arr_54),
    .io_arr_55(__m_fill_1_io_arr_55),
    .io_arr_56(__m_fill_1_io_arr_56),
    .io_arr_57(__m_fill_1_io_arr_57),
    .io_arr_58(__m_fill_1_io_arr_58),
    .io_arr_59(__m_fill_1_io_arr_59),
    .io_arr_60(__m_fill_1_io_arr_60),
    .io_arr_61(__m_fill_1_io_arr_61),
    .io_arr_62(__m_fill_1_io_arr_62),
    .io_arr_63(__m_fill_1_io_arr_63),
    .io_arr_64(__m_fill_1_io_arr_64),
    .io_arr_65(__m_fill_1_io_arr_65),
    .io_arr_66(__m_fill_1_io_arr_66),
    .io_arr_67(__m_fill_1_io_arr_67),
    .io_arr_68(__m_fill_1_io_arr_68),
    .io_arr_69(__m_fill_1_io_arr_69),
    .io_arr_70(__m_fill_1_io_arr_70),
    .io_arr_71(__m_fill_1_io_arr_71),
    .io_arr_72(__m_fill_1_io_arr_72),
    .io_arr_73(__m_fill_1_io_arr_73),
    .io_arr_74(__m_fill_1_io_arr_74),
    .io_arr_75(__m_fill_1_io_arr_75),
    .io_arr_76(__m_fill_1_io_arr_76),
    .io_arr_77(__m_fill_1_io_arr_77),
    .io_arr_78(__m_fill_1_io_arr_78),
    .io_arr_79(__m_fill_1_io_arr_79),
    .io_off(__m_fill_1_io_off),
    .io_valid(__m_fill_1_io_valid),
    .io_arr_out_0(__m_fill_1_io_arr_out_0),
    .io_arr_out_1(__m_fill_1_io_arr_out_1),
    .io_arr_out_2(__m_fill_1_io_arr_out_2),
    .io_arr_out_3(__m_fill_1_io_arr_out_3),
    .io_arr_out_4(__m_fill_1_io_arr_out_4),
    .io_arr_out_5(__m_fill_1_io_arr_out_5),
    .io_arr_out_6(__m_fill_1_io_arr_out_6),
    .io_arr_out_7(__m_fill_1_io_arr_out_7),
    .io_arr_out_8(__m_fill_1_io_arr_out_8),
    .io_arr_out_9(__m_fill_1_io_arr_out_9),
    .io_arr_out_10(__m_fill_1_io_arr_out_10),
    .io_arr_out_11(__m_fill_1_io_arr_out_11),
    .io_arr_out_12(__m_fill_1_io_arr_out_12),
    .io_arr_out_13(__m_fill_1_io_arr_out_13),
    .io_arr_out_14(__m_fill_1_io_arr_out_14),
    .io_arr_out_15(__m_fill_1_io_arr_out_15),
    .io_arr_out_16(__m_fill_1_io_arr_out_16),
    .io_arr_out_17(__m_fill_1_io_arr_out_17),
    .io_arr_out_18(__m_fill_1_io_arr_out_18),
    .io_arr_out_19(__m_fill_1_io_arr_out_19),
    .io_arr_out_20(__m_fill_1_io_arr_out_20),
    .io_arr_out_21(__m_fill_1_io_arr_out_21),
    .io_arr_out_22(__m_fill_1_io_arr_out_22),
    .io_arr_out_23(__m_fill_1_io_arr_out_23),
    .io_arr_out_24(__m_fill_1_io_arr_out_24),
    .io_arr_out_25(__m_fill_1_io_arr_out_25),
    .io_arr_out_26(__m_fill_1_io_arr_out_26),
    .io_arr_out_27(__m_fill_1_io_arr_out_27),
    .io_arr_out_28(__m_fill_1_io_arr_out_28),
    .io_arr_out_29(__m_fill_1_io_arr_out_29),
    .io_arr_out_30(__m_fill_1_io_arr_out_30),
    .io_arr_out_31(__m_fill_1_io_arr_out_31),
    .io_arr_out_32(__m_fill_1_io_arr_out_32),
    .io_arr_out_33(__m_fill_1_io_arr_out_33),
    .io_arr_out_34(__m_fill_1_io_arr_out_34),
    .io_arr_out_35(__m_fill_1_io_arr_out_35),
    .io_arr_out_36(__m_fill_1_io_arr_out_36),
    .io_arr_out_37(__m_fill_1_io_arr_out_37),
    .io_arr_out_38(__m_fill_1_io_arr_out_38),
    .io_arr_out_39(__m_fill_1_io_arr_out_39),
    .io_arr_out_40(__m_fill_1_io_arr_out_40),
    .io_arr_out_41(__m_fill_1_io_arr_out_41),
    .io_arr_out_42(__m_fill_1_io_arr_out_42),
    .io_arr_out_43(__m_fill_1_io_arr_out_43),
    .io_arr_out_44(__m_fill_1_io_arr_out_44),
    .io_arr_out_45(__m_fill_1_io_arr_out_45),
    .io_arr_out_46(__m_fill_1_io_arr_out_46),
    .io_arr_out_47(__m_fill_1_io_arr_out_47),
    .io_arr_out_48(__m_fill_1_io_arr_out_48),
    .io_arr_out_49(__m_fill_1_io_arr_out_49),
    .io_arr_out_50(__m_fill_1_io_arr_out_50),
    .io_arr_out_51(__m_fill_1_io_arr_out_51),
    .io_arr_out_52(__m_fill_1_io_arr_out_52),
    .io_arr_out_53(__m_fill_1_io_arr_out_53),
    .io_arr_out_54(__m_fill_1_io_arr_out_54),
    .io_arr_out_55(__m_fill_1_io_arr_out_55),
    .io_arr_out_56(__m_fill_1_io_arr_out_56),
    .io_arr_out_57(__m_fill_1_io_arr_out_57),
    .io_arr_out_58(__m_fill_1_io_arr_out_58),
    .io_arr_out_59(__m_fill_1_io_arr_out_59),
    .io_arr_out_60(__m_fill_1_io_arr_out_60),
    .io_arr_out_61(__m_fill_1_io_arr_out_61),
    .io_arr_out_62(__m_fill_1_io_arr_out_62),
    .io_arr_out_63(__m_fill_1_io_arr_out_63),
    .io_arr_out_64(__m_fill_1_io_arr_out_64),
    .io_arr_out_65(__m_fill_1_io_arr_out_65),
    .io_arr_out_66(__m_fill_1_io_arr_out_66),
    .io_arr_out_67(__m_fill_1_io_arr_out_67),
    .io_arr_out_68(__m_fill_1_io_arr_out_68),
    .io_arr_out_69(__m_fill_1_io_arr_out_69),
    .io_arr_out_70(__m_fill_1_io_arr_out_70),
    .io_arr_out_71(__m_fill_1_io_arr_out_71),
    .io_arr_out_72(__m_fill_1_io_arr_out_72),
    .io_arr_out_73(__m_fill_1_io_arr_out_73),
    .io_arr_out_74(__m_fill_1_io_arr_out_74),
    .io_arr_out_75(__m_fill_1_io_arr_out_75),
    .io_arr_out_76(__m_fill_1_io_arr_out_76),
    .io_arr_out_77(__m_fill_1_io_arr_out_77),
    .io_arr_out_78(__m_fill_1_io_arr_out_78),
    .io_arr_out_79(__m_fill_1_io_arr_out_79),
    .io_ready(__m_fill_1_io_ready)
  );
  fill __m_fill_2 ( // @[digest.scala 64:28]
    .clock(__m_fill_2_clock),
    .reset(__m_fill_2_reset),
    .io_value(__m_fill_2_io_value),
    .io_arr_0(__m_fill_2_io_arr_0),
    .io_arr_1(__m_fill_2_io_arr_1),
    .io_arr_2(__m_fill_2_io_arr_2),
    .io_arr_3(__m_fill_2_io_arr_3),
    .io_arr_4(__m_fill_2_io_arr_4),
    .io_arr_5(__m_fill_2_io_arr_5),
    .io_arr_6(__m_fill_2_io_arr_6),
    .io_arr_7(__m_fill_2_io_arr_7),
    .io_arr_8(__m_fill_2_io_arr_8),
    .io_arr_9(__m_fill_2_io_arr_9),
    .io_arr_10(__m_fill_2_io_arr_10),
    .io_arr_11(__m_fill_2_io_arr_11),
    .io_arr_12(__m_fill_2_io_arr_12),
    .io_arr_13(__m_fill_2_io_arr_13),
    .io_arr_14(__m_fill_2_io_arr_14),
    .io_arr_15(__m_fill_2_io_arr_15),
    .io_arr_16(__m_fill_2_io_arr_16),
    .io_arr_17(__m_fill_2_io_arr_17),
    .io_arr_18(__m_fill_2_io_arr_18),
    .io_arr_19(__m_fill_2_io_arr_19),
    .io_arr_20(__m_fill_2_io_arr_20),
    .io_arr_21(__m_fill_2_io_arr_21),
    .io_arr_22(__m_fill_2_io_arr_22),
    .io_arr_23(__m_fill_2_io_arr_23),
    .io_arr_24(__m_fill_2_io_arr_24),
    .io_arr_25(__m_fill_2_io_arr_25),
    .io_arr_26(__m_fill_2_io_arr_26),
    .io_arr_27(__m_fill_2_io_arr_27),
    .io_arr_28(__m_fill_2_io_arr_28),
    .io_arr_29(__m_fill_2_io_arr_29),
    .io_arr_30(__m_fill_2_io_arr_30),
    .io_arr_31(__m_fill_2_io_arr_31),
    .io_arr_32(__m_fill_2_io_arr_32),
    .io_arr_33(__m_fill_2_io_arr_33),
    .io_arr_34(__m_fill_2_io_arr_34),
    .io_arr_35(__m_fill_2_io_arr_35),
    .io_arr_36(__m_fill_2_io_arr_36),
    .io_arr_37(__m_fill_2_io_arr_37),
    .io_arr_38(__m_fill_2_io_arr_38),
    .io_arr_39(__m_fill_2_io_arr_39),
    .io_arr_40(__m_fill_2_io_arr_40),
    .io_arr_41(__m_fill_2_io_arr_41),
    .io_arr_42(__m_fill_2_io_arr_42),
    .io_arr_43(__m_fill_2_io_arr_43),
    .io_arr_44(__m_fill_2_io_arr_44),
    .io_arr_45(__m_fill_2_io_arr_45),
    .io_arr_46(__m_fill_2_io_arr_46),
    .io_arr_47(__m_fill_2_io_arr_47),
    .io_arr_48(__m_fill_2_io_arr_48),
    .io_arr_49(__m_fill_2_io_arr_49),
    .io_arr_50(__m_fill_2_io_arr_50),
    .io_arr_51(__m_fill_2_io_arr_51),
    .io_arr_52(__m_fill_2_io_arr_52),
    .io_arr_53(__m_fill_2_io_arr_53),
    .io_arr_54(__m_fill_2_io_arr_54),
    .io_arr_55(__m_fill_2_io_arr_55),
    .io_arr_56(__m_fill_2_io_arr_56),
    .io_arr_57(__m_fill_2_io_arr_57),
    .io_arr_58(__m_fill_2_io_arr_58),
    .io_arr_59(__m_fill_2_io_arr_59),
    .io_arr_60(__m_fill_2_io_arr_60),
    .io_arr_61(__m_fill_2_io_arr_61),
    .io_arr_62(__m_fill_2_io_arr_62),
    .io_arr_63(__m_fill_2_io_arr_63),
    .io_arr_64(__m_fill_2_io_arr_64),
    .io_arr_65(__m_fill_2_io_arr_65),
    .io_arr_66(__m_fill_2_io_arr_66),
    .io_arr_67(__m_fill_2_io_arr_67),
    .io_arr_68(__m_fill_2_io_arr_68),
    .io_arr_69(__m_fill_2_io_arr_69),
    .io_arr_70(__m_fill_2_io_arr_70),
    .io_arr_71(__m_fill_2_io_arr_71),
    .io_arr_72(__m_fill_2_io_arr_72),
    .io_arr_73(__m_fill_2_io_arr_73),
    .io_arr_74(__m_fill_2_io_arr_74),
    .io_arr_75(__m_fill_2_io_arr_75),
    .io_arr_76(__m_fill_2_io_arr_76),
    .io_arr_77(__m_fill_2_io_arr_77),
    .io_arr_78(__m_fill_2_io_arr_78),
    .io_arr_79(__m_fill_2_io_arr_79),
    .io_off(__m_fill_2_io_off),
    .io_valid(__m_fill_2_io_valid),
    .io_arr_out_0(__m_fill_2_io_arr_out_0),
    .io_arr_out_1(__m_fill_2_io_arr_out_1),
    .io_arr_out_2(__m_fill_2_io_arr_out_2),
    .io_arr_out_3(__m_fill_2_io_arr_out_3),
    .io_arr_out_4(__m_fill_2_io_arr_out_4),
    .io_arr_out_5(__m_fill_2_io_arr_out_5),
    .io_arr_out_6(__m_fill_2_io_arr_out_6),
    .io_arr_out_7(__m_fill_2_io_arr_out_7),
    .io_arr_out_8(__m_fill_2_io_arr_out_8),
    .io_arr_out_9(__m_fill_2_io_arr_out_9),
    .io_arr_out_10(__m_fill_2_io_arr_out_10),
    .io_arr_out_11(__m_fill_2_io_arr_out_11),
    .io_arr_out_12(__m_fill_2_io_arr_out_12),
    .io_arr_out_13(__m_fill_2_io_arr_out_13),
    .io_arr_out_14(__m_fill_2_io_arr_out_14),
    .io_arr_out_15(__m_fill_2_io_arr_out_15),
    .io_arr_out_16(__m_fill_2_io_arr_out_16),
    .io_arr_out_17(__m_fill_2_io_arr_out_17),
    .io_arr_out_18(__m_fill_2_io_arr_out_18),
    .io_arr_out_19(__m_fill_2_io_arr_out_19),
    .io_arr_out_20(__m_fill_2_io_arr_out_20),
    .io_arr_out_21(__m_fill_2_io_arr_out_21),
    .io_arr_out_22(__m_fill_2_io_arr_out_22),
    .io_arr_out_23(__m_fill_2_io_arr_out_23),
    .io_arr_out_24(__m_fill_2_io_arr_out_24),
    .io_arr_out_25(__m_fill_2_io_arr_out_25),
    .io_arr_out_26(__m_fill_2_io_arr_out_26),
    .io_arr_out_27(__m_fill_2_io_arr_out_27),
    .io_arr_out_28(__m_fill_2_io_arr_out_28),
    .io_arr_out_29(__m_fill_2_io_arr_out_29),
    .io_arr_out_30(__m_fill_2_io_arr_out_30),
    .io_arr_out_31(__m_fill_2_io_arr_out_31),
    .io_arr_out_32(__m_fill_2_io_arr_out_32),
    .io_arr_out_33(__m_fill_2_io_arr_out_33),
    .io_arr_out_34(__m_fill_2_io_arr_out_34),
    .io_arr_out_35(__m_fill_2_io_arr_out_35),
    .io_arr_out_36(__m_fill_2_io_arr_out_36),
    .io_arr_out_37(__m_fill_2_io_arr_out_37),
    .io_arr_out_38(__m_fill_2_io_arr_out_38),
    .io_arr_out_39(__m_fill_2_io_arr_out_39),
    .io_arr_out_40(__m_fill_2_io_arr_out_40),
    .io_arr_out_41(__m_fill_2_io_arr_out_41),
    .io_arr_out_42(__m_fill_2_io_arr_out_42),
    .io_arr_out_43(__m_fill_2_io_arr_out_43),
    .io_arr_out_44(__m_fill_2_io_arr_out_44),
    .io_arr_out_45(__m_fill_2_io_arr_out_45),
    .io_arr_out_46(__m_fill_2_io_arr_out_46),
    .io_arr_out_47(__m_fill_2_io_arr_out_47),
    .io_arr_out_48(__m_fill_2_io_arr_out_48),
    .io_arr_out_49(__m_fill_2_io_arr_out_49),
    .io_arr_out_50(__m_fill_2_io_arr_out_50),
    .io_arr_out_51(__m_fill_2_io_arr_out_51),
    .io_arr_out_52(__m_fill_2_io_arr_out_52),
    .io_arr_out_53(__m_fill_2_io_arr_out_53),
    .io_arr_out_54(__m_fill_2_io_arr_out_54),
    .io_arr_out_55(__m_fill_2_io_arr_out_55),
    .io_arr_out_56(__m_fill_2_io_arr_out_56),
    .io_arr_out_57(__m_fill_2_io_arr_out_57),
    .io_arr_out_58(__m_fill_2_io_arr_out_58),
    .io_arr_out_59(__m_fill_2_io_arr_out_59),
    .io_arr_out_60(__m_fill_2_io_arr_out_60),
    .io_arr_out_61(__m_fill_2_io_arr_out_61),
    .io_arr_out_62(__m_fill_2_io_arr_out_62),
    .io_arr_out_63(__m_fill_2_io_arr_out_63),
    .io_arr_out_64(__m_fill_2_io_arr_out_64),
    .io_arr_out_65(__m_fill_2_io_arr_out_65),
    .io_arr_out_66(__m_fill_2_io_arr_out_66),
    .io_arr_out_67(__m_fill_2_io_arr_out_67),
    .io_arr_out_68(__m_fill_2_io_arr_out_68),
    .io_arr_out_69(__m_fill_2_io_arr_out_69),
    .io_arr_out_70(__m_fill_2_io_arr_out_70),
    .io_arr_out_71(__m_fill_2_io_arr_out_71),
    .io_arr_out_72(__m_fill_2_io_arr_out_72),
    .io_arr_out_73(__m_fill_2_io_arr_out_73),
    .io_arr_out_74(__m_fill_2_io_arr_out_74),
    .io_arr_out_75(__m_fill_2_io_arr_out_75),
    .io_arr_out_76(__m_fill_2_io_arr_out_76),
    .io_arr_out_77(__m_fill_2_io_arr_out_77),
    .io_arr_out_78(__m_fill_2_io_arr_out_78),
    .io_arr_out_79(__m_fill_2_io_arr_out_79),
    .io_ready(__m_fill_2_io_ready)
  );
  fill __m_fill_3 ( // @[digest.scala 69:28]
    .clock(__m_fill_3_clock),
    .reset(__m_fill_3_reset),
    .io_value(__m_fill_3_io_value),
    .io_arr_0(__m_fill_3_io_arr_0),
    .io_arr_1(__m_fill_3_io_arr_1),
    .io_arr_2(__m_fill_3_io_arr_2),
    .io_arr_3(__m_fill_3_io_arr_3),
    .io_arr_4(__m_fill_3_io_arr_4),
    .io_arr_5(__m_fill_3_io_arr_5),
    .io_arr_6(__m_fill_3_io_arr_6),
    .io_arr_7(__m_fill_3_io_arr_7),
    .io_arr_8(__m_fill_3_io_arr_8),
    .io_arr_9(__m_fill_3_io_arr_9),
    .io_arr_10(__m_fill_3_io_arr_10),
    .io_arr_11(__m_fill_3_io_arr_11),
    .io_arr_12(__m_fill_3_io_arr_12),
    .io_arr_13(__m_fill_3_io_arr_13),
    .io_arr_14(__m_fill_3_io_arr_14),
    .io_arr_15(__m_fill_3_io_arr_15),
    .io_arr_16(__m_fill_3_io_arr_16),
    .io_arr_17(__m_fill_3_io_arr_17),
    .io_arr_18(__m_fill_3_io_arr_18),
    .io_arr_19(__m_fill_3_io_arr_19),
    .io_arr_20(__m_fill_3_io_arr_20),
    .io_arr_21(__m_fill_3_io_arr_21),
    .io_arr_22(__m_fill_3_io_arr_22),
    .io_arr_23(__m_fill_3_io_arr_23),
    .io_arr_24(__m_fill_3_io_arr_24),
    .io_arr_25(__m_fill_3_io_arr_25),
    .io_arr_26(__m_fill_3_io_arr_26),
    .io_arr_27(__m_fill_3_io_arr_27),
    .io_arr_28(__m_fill_3_io_arr_28),
    .io_arr_29(__m_fill_3_io_arr_29),
    .io_arr_30(__m_fill_3_io_arr_30),
    .io_arr_31(__m_fill_3_io_arr_31),
    .io_arr_32(__m_fill_3_io_arr_32),
    .io_arr_33(__m_fill_3_io_arr_33),
    .io_arr_34(__m_fill_3_io_arr_34),
    .io_arr_35(__m_fill_3_io_arr_35),
    .io_arr_36(__m_fill_3_io_arr_36),
    .io_arr_37(__m_fill_3_io_arr_37),
    .io_arr_38(__m_fill_3_io_arr_38),
    .io_arr_39(__m_fill_3_io_arr_39),
    .io_arr_40(__m_fill_3_io_arr_40),
    .io_arr_41(__m_fill_3_io_arr_41),
    .io_arr_42(__m_fill_3_io_arr_42),
    .io_arr_43(__m_fill_3_io_arr_43),
    .io_arr_44(__m_fill_3_io_arr_44),
    .io_arr_45(__m_fill_3_io_arr_45),
    .io_arr_46(__m_fill_3_io_arr_46),
    .io_arr_47(__m_fill_3_io_arr_47),
    .io_arr_48(__m_fill_3_io_arr_48),
    .io_arr_49(__m_fill_3_io_arr_49),
    .io_arr_50(__m_fill_3_io_arr_50),
    .io_arr_51(__m_fill_3_io_arr_51),
    .io_arr_52(__m_fill_3_io_arr_52),
    .io_arr_53(__m_fill_3_io_arr_53),
    .io_arr_54(__m_fill_3_io_arr_54),
    .io_arr_55(__m_fill_3_io_arr_55),
    .io_arr_56(__m_fill_3_io_arr_56),
    .io_arr_57(__m_fill_3_io_arr_57),
    .io_arr_58(__m_fill_3_io_arr_58),
    .io_arr_59(__m_fill_3_io_arr_59),
    .io_arr_60(__m_fill_3_io_arr_60),
    .io_arr_61(__m_fill_3_io_arr_61),
    .io_arr_62(__m_fill_3_io_arr_62),
    .io_arr_63(__m_fill_3_io_arr_63),
    .io_arr_64(__m_fill_3_io_arr_64),
    .io_arr_65(__m_fill_3_io_arr_65),
    .io_arr_66(__m_fill_3_io_arr_66),
    .io_arr_67(__m_fill_3_io_arr_67),
    .io_arr_68(__m_fill_3_io_arr_68),
    .io_arr_69(__m_fill_3_io_arr_69),
    .io_arr_70(__m_fill_3_io_arr_70),
    .io_arr_71(__m_fill_3_io_arr_71),
    .io_arr_72(__m_fill_3_io_arr_72),
    .io_arr_73(__m_fill_3_io_arr_73),
    .io_arr_74(__m_fill_3_io_arr_74),
    .io_arr_75(__m_fill_3_io_arr_75),
    .io_arr_76(__m_fill_3_io_arr_76),
    .io_arr_77(__m_fill_3_io_arr_77),
    .io_arr_78(__m_fill_3_io_arr_78),
    .io_arr_79(__m_fill_3_io_arr_79),
    .io_off(__m_fill_3_io_off),
    .io_valid(__m_fill_3_io_valid),
    .io_arr_out_0(__m_fill_3_io_arr_out_0),
    .io_arr_out_1(__m_fill_3_io_arr_out_1),
    .io_arr_out_2(__m_fill_3_io_arr_out_2),
    .io_arr_out_3(__m_fill_3_io_arr_out_3),
    .io_arr_out_4(__m_fill_3_io_arr_out_4),
    .io_arr_out_5(__m_fill_3_io_arr_out_5),
    .io_arr_out_6(__m_fill_3_io_arr_out_6),
    .io_arr_out_7(__m_fill_3_io_arr_out_7),
    .io_arr_out_8(__m_fill_3_io_arr_out_8),
    .io_arr_out_9(__m_fill_3_io_arr_out_9),
    .io_arr_out_10(__m_fill_3_io_arr_out_10),
    .io_arr_out_11(__m_fill_3_io_arr_out_11),
    .io_arr_out_12(__m_fill_3_io_arr_out_12),
    .io_arr_out_13(__m_fill_3_io_arr_out_13),
    .io_arr_out_14(__m_fill_3_io_arr_out_14),
    .io_arr_out_15(__m_fill_3_io_arr_out_15),
    .io_arr_out_16(__m_fill_3_io_arr_out_16),
    .io_arr_out_17(__m_fill_3_io_arr_out_17),
    .io_arr_out_18(__m_fill_3_io_arr_out_18),
    .io_arr_out_19(__m_fill_3_io_arr_out_19),
    .io_arr_out_20(__m_fill_3_io_arr_out_20),
    .io_arr_out_21(__m_fill_3_io_arr_out_21),
    .io_arr_out_22(__m_fill_3_io_arr_out_22),
    .io_arr_out_23(__m_fill_3_io_arr_out_23),
    .io_arr_out_24(__m_fill_3_io_arr_out_24),
    .io_arr_out_25(__m_fill_3_io_arr_out_25),
    .io_arr_out_26(__m_fill_3_io_arr_out_26),
    .io_arr_out_27(__m_fill_3_io_arr_out_27),
    .io_arr_out_28(__m_fill_3_io_arr_out_28),
    .io_arr_out_29(__m_fill_3_io_arr_out_29),
    .io_arr_out_30(__m_fill_3_io_arr_out_30),
    .io_arr_out_31(__m_fill_3_io_arr_out_31),
    .io_arr_out_32(__m_fill_3_io_arr_out_32),
    .io_arr_out_33(__m_fill_3_io_arr_out_33),
    .io_arr_out_34(__m_fill_3_io_arr_out_34),
    .io_arr_out_35(__m_fill_3_io_arr_out_35),
    .io_arr_out_36(__m_fill_3_io_arr_out_36),
    .io_arr_out_37(__m_fill_3_io_arr_out_37),
    .io_arr_out_38(__m_fill_3_io_arr_out_38),
    .io_arr_out_39(__m_fill_3_io_arr_out_39),
    .io_arr_out_40(__m_fill_3_io_arr_out_40),
    .io_arr_out_41(__m_fill_3_io_arr_out_41),
    .io_arr_out_42(__m_fill_3_io_arr_out_42),
    .io_arr_out_43(__m_fill_3_io_arr_out_43),
    .io_arr_out_44(__m_fill_3_io_arr_out_44),
    .io_arr_out_45(__m_fill_3_io_arr_out_45),
    .io_arr_out_46(__m_fill_3_io_arr_out_46),
    .io_arr_out_47(__m_fill_3_io_arr_out_47),
    .io_arr_out_48(__m_fill_3_io_arr_out_48),
    .io_arr_out_49(__m_fill_3_io_arr_out_49),
    .io_arr_out_50(__m_fill_3_io_arr_out_50),
    .io_arr_out_51(__m_fill_3_io_arr_out_51),
    .io_arr_out_52(__m_fill_3_io_arr_out_52),
    .io_arr_out_53(__m_fill_3_io_arr_out_53),
    .io_arr_out_54(__m_fill_3_io_arr_out_54),
    .io_arr_out_55(__m_fill_3_io_arr_out_55),
    .io_arr_out_56(__m_fill_3_io_arr_out_56),
    .io_arr_out_57(__m_fill_3_io_arr_out_57),
    .io_arr_out_58(__m_fill_3_io_arr_out_58),
    .io_arr_out_59(__m_fill_3_io_arr_out_59),
    .io_arr_out_60(__m_fill_3_io_arr_out_60),
    .io_arr_out_61(__m_fill_3_io_arr_out_61),
    .io_arr_out_62(__m_fill_3_io_arr_out_62),
    .io_arr_out_63(__m_fill_3_io_arr_out_63),
    .io_arr_out_64(__m_fill_3_io_arr_out_64),
    .io_arr_out_65(__m_fill_3_io_arr_out_65),
    .io_arr_out_66(__m_fill_3_io_arr_out_66),
    .io_arr_out_67(__m_fill_3_io_arr_out_67),
    .io_arr_out_68(__m_fill_3_io_arr_out_68),
    .io_arr_out_69(__m_fill_3_io_arr_out_69),
    .io_arr_out_70(__m_fill_3_io_arr_out_70),
    .io_arr_out_71(__m_fill_3_io_arr_out_71),
    .io_arr_out_72(__m_fill_3_io_arr_out_72),
    .io_arr_out_73(__m_fill_3_io_arr_out_73),
    .io_arr_out_74(__m_fill_3_io_arr_out_74),
    .io_arr_out_75(__m_fill_3_io_arr_out_75),
    .io_arr_out_76(__m_fill_3_io_arr_out_76),
    .io_arr_out_77(__m_fill_3_io_arr_out_77),
    .io_arr_out_78(__m_fill_3_io_arr_out_78),
    .io_arr_out_79(__m_fill_3_io_arr_out_79),
    .io_ready(__m_fill_3_io_ready)
  );
  fill __m_fill_4 ( // @[digest.scala 74:28]
    .clock(__m_fill_4_clock),
    .reset(__m_fill_4_reset),
    .io_value(__m_fill_4_io_value),
    .io_arr_0(__m_fill_4_io_arr_0),
    .io_arr_1(__m_fill_4_io_arr_1),
    .io_arr_2(__m_fill_4_io_arr_2),
    .io_arr_3(__m_fill_4_io_arr_3),
    .io_arr_4(__m_fill_4_io_arr_4),
    .io_arr_5(__m_fill_4_io_arr_5),
    .io_arr_6(__m_fill_4_io_arr_6),
    .io_arr_7(__m_fill_4_io_arr_7),
    .io_arr_8(__m_fill_4_io_arr_8),
    .io_arr_9(__m_fill_4_io_arr_9),
    .io_arr_10(__m_fill_4_io_arr_10),
    .io_arr_11(__m_fill_4_io_arr_11),
    .io_arr_12(__m_fill_4_io_arr_12),
    .io_arr_13(__m_fill_4_io_arr_13),
    .io_arr_14(__m_fill_4_io_arr_14),
    .io_arr_15(__m_fill_4_io_arr_15),
    .io_arr_16(__m_fill_4_io_arr_16),
    .io_arr_17(__m_fill_4_io_arr_17),
    .io_arr_18(__m_fill_4_io_arr_18),
    .io_arr_19(__m_fill_4_io_arr_19),
    .io_arr_20(__m_fill_4_io_arr_20),
    .io_arr_21(__m_fill_4_io_arr_21),
    .io_arr_22(__m_fill_4_io_arr_22),
    .io_arr_23(__m_fill_4_io_arr_23),
    .io_arr_24(__m_fill_4_io_arr_24),
    .io_arr_25(__m_fill_4_io_arr_25),
    .io_arr_26(__m_fill_4_io_arr_26),
    .io_arr_27(__m_fill_4_io_arr_27),
    .io_arr_28(__m_fill_4_io_arr_28),
    .io_arr_29(__m_fill_4_io_arr_29),
    .io_arr_30(__m_fill_4_io_arr_30),
    .io_arr_31(__m_fill_4_io_arr_31),
    .io_arr_32(__m_fill_4_io_arr_32),
    .io_arr_33(__m_fill_4_io_arr_33),
    .io_arr_34(__m_fill_4_io_arr_34),
    .io_arr_35(__m_fill_4_io_arr_35),
    .io_arr_36(__m_fill_4_io_arr_36),
    .io_arr_37(__m_fill_4_io_arr_37),
    .io_arr_38(__m_fill_4_io_arr_38),
    .io_arr_39(__m_fill_4_io_arr_39),
    .io_arr_40(__m_fill_4_io_arr_40),
    .io_arr_41(__m_fill_4_io_arr_41),
    .io_arr_42(__m_fill_4_io_arr_42),
    .io_arr_43(__m_fill_4_io_arr_43),
    .io_arr_44(__m_fill_4_io_arr_44),
    .io_arr_45(__m_fill_4_io_arr_45),
    .io_arr_46(__m_fill_4_io_arr_46),
    .io_arr_47(__m_fill_4_io_arr_47),
    .io_arr_48(__m_fill_4_io_arr_48),
    .io_arr_49(__m_fill_4_io_arr_49),
    .io_arr_50(__m_fill_4_io_arr_50),
    .io_arr_51(__m_fill_4_io_arr_51),
    .io_arr_52(__m_fill_4_io_arr_52),
    .io_arr_53(__m_fill_4_io_arr_53),
    .io_arr_54(__m_fill_4_io_arr_54),
    .io_arr_55(__m_fill_4_io_arr_55),
    .io_arr_56(__m_fill_4_io_arr_56),
    .io_arr_57(__m_fill_4_io_arr_57),
    .io_arr_58(__m_fill_4_io_arr_58),
    .io_arr_59(__m_fill_4_io_arr_59),
    .io_arr_60(__m_fill_4_io_arr_60),
    .io_arr_61(__m_fill_4_io_arr_61),
    .io_arr_62(__m_fill_4_io_arr_62),
    .io_arr_63(__m_fill_4_io_arr_63),
    .io_arr_64(__m_fill_4_io_arr_64),
    .io_arr_65(__m_fill_4_io_arr_65),
    .io_arr_66(__m_fill_4_io_arr_66),
    .io_arr_67(__m_fill_4_io_arr_67),
    .io_arr_68(__m_fill_4_io_arr_68),
    .io_arr_69(__m_fill_4_io_arr_69),
    .io_arr_70(__m_fill_4_io_arr_70),
    .io_arr_71(__m_fill_4_io_arr_71),
    .io_arr_72(__m_fill_4_io_arr_72),
    .io_arr_73(__m_fill_4_io_arr_73),
    .io_arr_74(__m_fill_4_io_arr_74),
    .io_arr_75(__m_fill_4_io_arr_75),
    .io_arr_76(__m_fill_4_io_arr_76),
    .io_arr_77(__m_fill_4_io_arr_77),
    .io_arr_78(__m_fill_4_io_arr_78),
    .io_arr_79(__m_fill_4_io_arr_79),
    .io_off(__m_fill_4_io_off),
    .io_valid(__m_fill_4_io_valid),
    .io_arr_out_0(__m_fill_4_io_arr_out_0),
    .io_arr_out_1(__m_fill_4_io_arr_out_1),
    .io_arr_out_2(__m_fill_4_io_arr_out_2),
    .io_arr_out_3(__m_fill_4_io_arr_out_3),
    .io_arr_out_4(__m_fill_4_io_arr_out_4),
    .io_arr_out_5(__m_fill_4_io_arr_out_5),
    .io_arr_out_6(__m_fill_4_io_arr_out_6),
    .io_arr_out_7(__m_fill_4_io_arr_out_7),
    .io_arr_out_8(__m_fill_4_io_arr_out_8),
    .io_arr_out_9(__m_fill_4_io_arr_out_9),
    .io_arr_out_10(__m_fill_4_io_arr_out_10),
    .io_arr_out_11(__m_fill_4_io_arr_out_11),
    .io_arr_out_12(__m_fill_4_io_arr_out_12),
    .io_arr_out_13(__m_fill_4_io_arr_out_13),
    .io_arr_out_14(__m_fill_4_io_arr_out_14),
    .io_arr_out_15(__m_fill_4_io_arr_out_15),
    .io_arr_out_16(__m_fill_4_io_arr_out_16),
    .io_arr_out_17(__m_fill_4_io_arr_out_17),
    .io_arr_out_18(__m_fill_4_io_arr_out_18),
    .io_arr_out_19(__m_fill_4_io_arr_out_19),
    .io_arr_out_20(__m_fill_4_io_arr_out_20),
    .io_arr_out_21(__m_fill_4_io_arr_out_21),
    .io_arr_out_22(__m_fill_4_io_arr_out_22),
    .io_arr_out_23(__m_fill_4_io_arr_out_23),
    .io_arr_out_24(__m_fill_4_io_arr_out_24),
    .io_arr_out_25(__m_fill_4_io_arr_out_25),
    .io_arr_out_26(__m_fill_4_io_arr_out_26),
    .io_arr_out_27(__m_fill_4_io_arr_out_27),
    .io_arr_out_28(__m_fill_4_io_arr_out_28),
    .io_arr_out_29(__m_fill_4_io_arr_out_29),
    .io_arr_out_30(__m_fill_4_io_arr_out_30),
    .io_arr_out_31(__m_fill_4_io_arr_out_31),
    .io_arr_out_32(__m_fill_4_io_arr_out_32),
    .io_arr_out_33(__m_fill_4_io_arr_out_33),
    .io_arr_out_34(__m_fill_4_io_arr_out_34),
    .io_arr_out_35(__m_fill_4_io_arr_out_35),
    .io_arr_out_36(__m_fill_4_io_arr_out_36),
    .io_arr_out_37(__m_fill_4_io_arr_out_37),
    .io_arr_out_38(__m_fill_4_io_arr_out_38),
    .io_arr_out_39(__m_fill_4_io_arr_out_39),
    .io_arr_out_40(__m_fill_4_io_arr_out_40),
    .io_arr_out_41(__m_fill_4_io_arr_out_41),
    .io_arr_out_42(__m_fill_4_io_arr_out_42),
    .io_arr_out_43(__m_fill_4_io_arr_out_43),
    .io_arr_out_44(__m_fill_4_io_arr_out_44),
    .io_arr_out_45(__m_fill_4_io_arr_out_45),
    .io_arr_out_46(__m_fill_4_io_arr_out_46),
    .io_arr_out_47(__m_fill_4_io_arr_out_47),
    .io_arr_out_48(__m_fill_4_io_arr_out_48),
    .io_arr_out_49(__m_fill_4_io_arr_out_49),
    .io_arr_out_50(__m_fill_4_io_arr_out_50),
    .io_arr_out_51(__m_fill_4_io_arr_out_51),
    .io_arr_out_52(__m_fill_4_io_arr_out_52),
    .io_arr_out_53(__m_fill_4_io_arr_out_53),
    .io_arr_out_54(__m_fill_4_io_arr_out_54),
    .io_arr_out_55(__m_fill_4_io_arr_out_55),
    .io_arr_out_56(__m_fill_4_io_arr_out_56),
    .io_arr_out_57(__m_fill_4_io_arr_out_57),
    .io_arr_out_58(__m_fill_4_io_arr_out_58),
    .io_arr_out_59(__m_fill_4_io_arr_out_59),
    .io_arr_out_60(__m_fill_4_io_arr_out_60),
    .io_arr_out_61(__m_fill_4_io_arr_out_61),
    .io_arr_out_62(__m_fill_4_io_arr_out_62),
    .io_arr_out_63(__m_fill_4_io_arr_out_63),
    .io_arr_out_64(__m_fill_4_io_arr_out_64),
    .io_arr_out_65(__m_fill_4_io_arr_out_65),
    .io_arr_out_66(__m_fill_4_io_arr_out_66),
    .io_arr_out_67(__m_fill_4_io_arr_out_67),
    .io_arr_out_68(__m_fill_4_io_arr_out_68),
    .io_arr_out_69(__m_fill_4_io_arr_out_69),
    .io_arr_out_70(__m_fill_4_io_arr_out_70),
    .io_arr_out_71(__m_fill_4_io_arr_out_71),
    .io_arr_out_72(__m_fill_4_io_arr_out_72),
    .io_arr_out_73(__m_fill_4_io_arr_out_73),
    .io_arr_out_74(__m_fill_4_io_arr_out_74),
    .io_arr_out_75(__m_fill_4_io_arr_out_75),
    .io_arr_out_76(__m_fill_4_io_arr_out_76),
    .io_arr_out_77(__m_fill_4_io_arr_out_77),
    .io_arr_out_78(__m_fill_4_io_arr_out_78),
    .io_arr_out_79(__m_fill_4_io_arr_out_79),
    .io_ready(__m_fill_4_io_ready)
  );
  assign io_bytes_out_0 = bytes_0; // @[digest.scala 22:18]
  assign io_bytes_out_1 = bytes_1; // @[digest.scala 22:18]
  assign io_bytes_out_2 = bytes_2; // @[digest.scala 22:18]
  assign io_bytes_out_3 = bytes_3; // @[digest.scala 22:18]
  assign io_bytes_out_4 = bytes_4; // @[digest.scala 22:18]
  assign io_bytes_out_5 = bytes_5; // @[digest.scala 22:18]
  assign io_bytes_out_6 = bytes_6; // @[digest.scala 22:18]
  assign io_bytes_out_7 = bytes_7; // @[digest.scala 22:18]
  assign io_bytes_out_8 = bytes_8; // @[digest.scala 22:18]
  assign io_bytes_out_9 = bytes_9; // @[digest.scala 22:18]
  assign io_bytes_out_10 = bytes_10; // @[digest.scala 22:18]
  assign io_bytes_out_11 = bytes_11; // @[digest.scala 22:18]
  assign io_bytes_out_12 = bytes_12; // @[digest.scala 22:18]
  assign io_bytes_out_13 = bytes_13; // @[digest.scala 22:18]
  assign io_bytes_out_14 = bytes_14; // @[digest.scala 22:18]
  assign io_bytes_out_15 = bytes_15; // @[digest.scala 22:18]
  assign io_bytes_out_16 = bytes_16; // @[digest.scala 22:18]
  assign io_bytes_out_17 = bytes_17; // @[digest.scala 22:18]
  assign io_bytes_out_18 = bytes_18; // @[digest.scala 22:18]
  assign io_bytes_out_19 = bytes_19; // @[digest.scala 22:18]
  assign io_bytes_out_20 = bytes_20; // @[digest.scala 22:18]
  assign io_bytes_out_21 = bytes_21; // @[digest.scala 22:18]
  assign io_bytes_out_22 = bytes_22; // @[digest.scala 22:18]
  assign io_bytes_out_23 = bytes_23; // @[digest.scala 22:18]
  assign io_bytes_out_24 = bytes_24; // @[digest.scala 22:18]
  assign io_bytes_out_25 = bytes_25; // @[digest.scala 22:18]
  assign io_bytes_out_26 = bytes_26; // @[digest.scala 22:18]
  assign io_bytes_out_27 = bytes_27; // @[digest.scala 22:18]
  assign io_bytes_out_28 = bytes_28; // @[digest.scala 22:18]
  assign io_bytes_out_29 = bytes_29; // @[digest.scala 22:18]
  assign io_bytes_out_30 = bytes_30; // @[digest.scala 22:18]
  assign io_bytes_out_31 = bytes_31; // @[digest.scala 22:18]
  assign io_bytes_out_32 = bytes_32; // @[digest.scala 22:18]
  assign io_bytes_out_33 = bytes_33; // @[digest.scala 22:18]
  assign io_bytes_out_34 = bytes_34; // @[digest.scala 22:18]
  assign io_bytes_out_35 = bytes_35; // @[digest.scala 22:18]
  assign io_bytes_out_36 = bytes_36; // @[digest.scala 22:18]
  assign io_bytes_out_37 = bytes_37; // @[digest.scala 22:18]
  assign io_bytes_out_38 = bytes_38; // @[digest.scala 22:18]
  assign io_bytes_out_39 = bytes_39; // @[digest.scala 22:18]
  assign io_bytes_out_40 = bytes_40; // @[digest.scala 22:18]
  assign io_bytes_out_41 = bytes_41; // @[digest.scala 22:18]
  assign io_bytes_out_42 = bytes_42; // @[digest.scala 22:18]
  assign io_bytes_out_43 = bytes_43; // @[digest.scala 22:18]
  assign io_bytes_out_44 = bytes_44; // @[digest.scala 22:18]
  assign io_bytes_out_45 = bytes_45; // @[digest.scala 22:18]
  assign io_bytes_out_46 = bytes_46; // @[digest.scala 22:18]
  assign io_bytes_out_47 = bytes_47; // @[digest.scala 22:18]
  assign io_bytes_out_48 = bytes_48; // @[digest.scala 22:18]
  assign io_bytes_out_49 = bytes_49; // @[digest.scala 22:18]
  assign io_bytes_out_50 = bytes_50; // @[digest.scala 22:18]
  assign io_bytes_out_51 = bytes_51; // @[digest.scala 22:18]
  assign io_bytes_out_52 = bytes_52; // @[digest.scala 22:18]
  assign io_bytes_out_53 = bytes_53; // @[digest.scala 22:18]
  assign io_bytes_out_54 = bytes_54; // @[digest.scala 22:18]
  assign io_bytes_out_55 = bytes_55; // @[digest.scala 22:18]
  assign io_bytes_out_56 = bytes_56; // @[digest.scala 22:18]
  assign io_bytes_out_57 = bytes_57; // @[digest.scala 22:18]
  assign io_bytes_out_58 = bytes_58; // @[digest.scala 22:18]
  assign io_bytes_out_59 = bytes_59; // @[digest.scala 22:18]
  assign io_bytes_out_60 = bytes_60; // @[digest.scala 22:18]
  assign io_bytes_out_61 = bytes_61; // @[digest.scala 22:18]
  assign io_bytes_out_62 = bytes_62; // @[digest.scala 22:18]
  assign io_bytes_out_63 = bytes_63; // @[digest.scala 22:18]
  assign io_bytes_out_64 = bytes_64; // @[digest.scala 22:18]
  assign io_bytes_out_65 = bytes_65; // @[digest.scala 22:18]
  assign io_bytes_out_66 = bytes_66; // @[digest.scala 22:18]
  assign io_bytes_out_67 = bytes_67; // @[digest.scala 22:18]
  assign io_bytes_out_68 = bytes_68; // @[digest.scala 22:18]
  assign io_bytes_out_69 = bytes_69; // @[digest.scala 22:18]
  assign io_bytes_out_70 = bytes_70; // @[digest.scala 22:18]
  assign io_bytes_out_71 = bytes_71; // @[digest.scala 22:18]
  assign io_bytes_out_72 = bytes_72; // @[digest.scala 22:18]
  assign io_bytes_out_73 = bytes_73; // @[digest.scala 22:18]
  assign io_bytes_out_74 = bytes_74; // @[digest.scala 22:18]
  assign io_bytes_out_75 = bytes_75; // @[digest.scala 22:18]
  assign io_bytes_out_76 = bytes_76; // @[digest.scala 22:18]
  assign io_bytes_out_77 = bytes_77; // @[digest.scala 22:18]
  assign io_bytes_out_78 = bytes_78; // @[digest.scala 22:18]
  assign io_bytes_out_79 = bytes_79; // @[digest.scala 22:18]
  assign io_ready = state == 6'h3b; // @[digest.scala 358:23]
  assign io_out_digest_0 = digest_0; // @[digest.scala 79:12]
  assign io_out_digest_1 = digest_1; // @[digest.scala 79:12]
  assign io_out_digest_2 = digest_2; // @[digest.scala 79:12]
  assign io_out_digest_3 = digest_3; // @[digest.scala 79:12]
  assign io_out_digest_4 = digest_4; // @[digest.scala 79:12]
  assign io_out_digest_5 = digest_5; // @[digest.scala 79:12]
  assign io_out_digest_6 = digest_6; // @[digest.scala 79:12]
  assign io_out_digest_7 = digest_7; // @[digest.scala 79:12]
  assign io_out_digest_8 = digest_8; // @[digest.scala 79:12]
  assign io_out_digest_9 = digest_9; // @[digest.scala 79:12]
  assign io_out_digest_10 = digest_10; // @[digest.scala 79:12]
  assign io_out_digest_11 = digest_11; // @[digest.scala 79:12]
  assign io_out_digest_12 = digest_12; // @[digest.scala 79:12]
  assign io_out_digest_13 = digest_13; // @[digest.scala 79:12]
  assign io_out_digest_14 = digest_14; // @[digest.scala 79:12]
  assign io_out_digest_15 = digest_15; // @[digest.scala 79:12]
  assign io_out_digest_16 = digest_16; // @[digest.scala 79:12]
  assign io_out_digest_17 = digest_17; // @[digest.scala 79:12]
  assign io_out_digest_18 = digest_18; // @[digest.scala 79:12]
  assign io_out_digest_19 = digest_19; // @[digest.scala 79:12]
  assign io_out_digest_20 = digest_20; // @[digest.scala 79:12]
  assign io_out_digest_21 = digest_21; // @[digest.scala 79:12]
  assign io_out_digest_22 = digest_22; // @[digest.scala 79:12]
  assign io_out_digest_23 = digest_23; // @[digest.scala 79:12]
  assign io_out_digest_24 = digest_24; // @[digest.scala 79:12]
  assign io_out_digest_25 = digest_25; // @[digest.scala 79:12]
  assign io_out_digest_26 = digest_26; // @[digest.scala 79:12]
  assign io_out_digest_27 = digest_27; // @[digest.scala 79:12]
  assign io_out_digest_28 = digest_28; // @[digest.scala 79:12]
  assign io_out_digest_29 = digest_29; // @[digest.scala 79:12]
  assign io_out_digest_30 = digest_30; // @[digest.scala 79:12]
  assign io_out_digest_31 = digest_31; // @[digest.scala 79:12]
  assign io_out_digest_32 = digest_32; // @[digest.scala 79:12]
  assign io_out_digest_33 = digest_33; // @[digest.scala 79:12]
  assign io_out_digest_34 = digest_34; // @[digest.scala 79:12]
  assign io_out_digest_35 = digest_35; // @[digest.scala 79:12]
  assign io_out_digest_36 = digest_36; // @[digest.scala 79:12]
  assign io_out_digest_37 = digest_37; // @[digest.scala 79:12]
  assign io_out_digest_38 = digest_38; // @[digest.scala 79:12]
  assign io_out_digest_39 = digest_39; // @[digest.scala 79:12]
  assign io_out_digest_40 = digest_40; // @[digest.scala 79:12]
  assign io_out_digest_41 = digest_41; // @[digest.scala 79:12]
  assign io_out_digest_42 = digest_42; // @[digest.scala 79:12]
  assign io_out_digest_43 = digest_43; // @[digest.scala 79:12]
  assign io_out_digest_44 = digest_44; // @[digest.scala 79:12]
  assign io_out_digest_45 = digest_45; // @[digest.scala 79:12]
  assign io_out_digest_46 = digest_46; // @[digest.scala 79:12]
  assign io_out_digest_47 = digest_47; // @[digest.scala 79:12]
  assign io_out_digest_48 = digest_48; // @[digest.scala 79:12]
  assign io_out_digest_49 = digest_49; // @[digest.scala 79:12]
  assign io_out_digest_50 = digest_50; // @[digest.scala 79:12]
  assign io_out_digest_51 = digest_51; // @[digest.scala 79:12]
  assign io_out_digest_52 = digest_52; // @[digest.scala 79:12]
  assign io_out_digest_53 = digest_53; // @[digest.scala 79:12]
  assign io_out_digest_54 = digest_54; // @[digest.scala 79:12]
  assign io_out_digest_55 = digest_55; // @[digest.scala 79:12]
  assign io_out_digest_56 = digest_56; // @[digest.scala 79:12]
  assign io_out_digest_57 = digest_57; // @[digest.scala 79:12]
  assign io_out_digest_58 = digest_58; // @[digest.scala 79:12]
  assign io_out_digest_59 = digest_59; // @[digest.scala 79:12]
  assign io_out_digest_60 = digest_60; // @[digest.scala 79:12]
  assign io_out_digest_61 = digest_61; // @[digest.scala 79:12]
  assign io_out_digest_62 = digest_62; // @[digest.scala 79:12]
  assign io_out_digest_63 = digest_63; // @[digest.scala 79:12]
  assign io_out_digest_64 = digest_64; // @[digest.scala 79:12]
  assign io_out_digest_65 = digest_65; // @[digest.scala 79:12]
  assign io_out_digest_66 = digest_66; // @[digest.scala 79:12]
  assign io_out_digest_67 = digest_67; // @[digest.scala 79:12]
  assign io_out_digest_68 = digest_68; // @[digest.scala 79:12]
  assign io_out_digest_69 = digest_69; // @[digest.scala 79:12]
  assign io_out_digest_70 = digest_70; // @[digest.scala 79:12]
  assign io_out_digest_71 = digest_71; // @[digest.scala 79:12]
  assign io_out_digest_72 = digest_72; // @[digest.scala 79:12]
  assign io_out_digest_73 = digest_73; // @[digest.scala 79:12]
  assign io_out_digest_74 = digest_74; // @[digest.scala 79:12]
  assign io_out_digest_75 = digest_75; // @[digest.scala 79:12]
  assign io_out_digest_76 = digest_76; // @[digest.scala 79:12]
  assign io_out_digest_77 = digest_77; // @[digest.scala 79:12]
  assign io_out_digest_78 = digest_78; // @[digest.scala 79:12]
  assign io_out_digest_79 = digest_79; // @[digest.scala 79:12]
  assign __m_rol_0_clock = clock;
  assign __m_rol_0_reset = reset;
  assign __m_rol_0_io_num = temp; // @[digest.scala 81:19 192:30]
  assign __m_rol_0_io_cnt = 32'sh1; // @[digest.scala 81:19 193:30]
  assign __m_rol_0_io_valid = 6'h3f == state ? 1'h0 : _GEN_33455; // @[digest.scala 81:19 44:24]
  assign __m_rol_1_clock = clock;
  assign __m_rol_1_reset = reset;
  assign __m_rol_1_io_num = a; // @[digest.scala 81:19 244:30]
  assign __m_rol_1_io_cnt = 32'sh5; // @[digest.scala 81:19 245:30]
  assign __m_rol_1_io_valid = 6'h3f == state ? 1'h0 : _GEN_33459; // @[digest.scala 81:19 48:24]
  assign __m_rol_2_clock = clock;
  assign __m_rol_2_reset = reset;
  assign __m_rol_2_io_num = b; // @[digest.scala 81:19 263:30]
  assign __m_rol_2_io_cnt = 32'sh1e; // @[digest.scala 81:19 264:30]
  assign __m_rol_2_io_valid = 6'h3f == state ? 1'h0 : _GEN_33462; // @[digest.scala 81:19 52:24]
  assign __m_fill_0_clock = clock;
  assign __m_fill_0_reset = reset;
  assign __m_fill_0_io_value = a; // @[digest.scala 81:19 304:33]
  assign __m_fill_0_io_arr_0 = digest_0; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_1 = digest_1; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_2 = digest_2; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_3 = digest_3; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_4 = digest_4; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_5 = digest_5; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_6 = digest_6; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_7 = digest_7; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_8 = digest_8; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_9 = digest_9; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_10 = digest_10; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_11 = digest_11; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_12 = digest_12; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_13 = digest_13; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_14 = digest_14; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_15 = digest_15; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_16 = digest_16; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_17 = digest_17; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_18 = digest_18; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_19 = digest_19; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_20 = digest_20; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_21 = digest_21; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_22 = digest_22; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_23 = digest_23; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_24 = digest_24; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_25 = digest_25; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_26 = digest_26; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_27 = digest_27; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_28 = digest_28; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_29 = digest_29; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_30 = digest_30; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_31 = digest_31; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_32 = digest_32; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_33 = digest_33; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_34 = digest_34; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_35 = digest_35; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_36 = digest_36; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_37 = digest_37; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_38 = digest_38; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_39 = digest_39; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_40 = digest_40; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_41 = digest_41; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_42 = digest_42; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_43 = digest_43; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_44 = digest_44; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_45 = digest_45; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_46 = digest_46; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_47 = digest_47; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_48 = digest_48; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_49 = digest_49; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_50 = digest_50; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_51 = digest_51; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_52 = digest_52; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_53 = digest_53; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_54 = digest_54; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_55 = digest_55; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_56 = digest_56; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_57 = digest_57; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_58 = digest_58; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_59 = digest_59; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_60 = digest_60; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_61 = digest_61; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_62 = digest_62; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_63 = digest_63; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_64 = digest_64; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_65 = digest_65; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_66 = digest_66; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_67 = digest_67; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_68 = digest_68; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_69 = digest_69; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_70 = digest_70; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_71 = digest_71; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_72 = digest_72; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_73 = digest_73; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_74 = digest_74; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_75 = digest_75; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_76 = digest_76; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_77 = digest_77; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_78 = digest_78; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_arr_79 = digest_79; // @[digest.scala 81:19 305:31]
  assign __m_fill_0_io_off = 32'sh0; // @[digest.scala 81:19 309:31]
  assign __m_fill_0_io_valid = 6'h3f == state ? 1'h0 : _GEN_33627; // @[digest.scala 81:19 58:25]
  assign __m_fill_1_clock = clock;
  assign __m_fill_1_reset = reset;
  assign __m_fill_1_io_value = b; // @[digest.scala 81:19 314:33]
  assign __m_fill_1_io_arr_0 = digest_0; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_1 = digest_1; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_2 = digest_2; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_3 = digest_3; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_4 = digest_4; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_5 = digest_5; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_6 = digest_6; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_7 = digest_7; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_8 = digest_8; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_9 = digest_9; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_10 = digest_10; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_11 = digest_11; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_12 = digest_12; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_13 = digest_13; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_14 = digest_14; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_15 = digest_15; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_16 = digest_16; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_17 = digest_17; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_18 = digest_18; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_19 = digest_19; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_20 = digest_20; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_21 = digest_21; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_22 = digest_22; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_23 = digest_23; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_24 = digest_24; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_25 = digest_25; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_26 = digest_26; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_27 = digest_27; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_28 = digest_28; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_29 = digest_29; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_30 = digest_30; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_31 = digest_31; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_32 = digest_32; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_33 = digest_33; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_34 = digest_34; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_35 = digest_35; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_36 = digest_36; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_37 = digest_37; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_38 = digest_38; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_39 = digest_39; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_40 = digest_40; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_41 = digest_41; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_42 = digest_42; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_43 = digest_43; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_44 = digest_44; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_45 = digest_45; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_46 = digest_46; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_47 = digest_47; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_48 = digest_48; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_49 = digest_49; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_50 = digest_50; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_51 = digest_51; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_52 = digest_52; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_53 = digest_53; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_54 = digest_54; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_55 = digest_55; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_56 = digest_56; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_57 = digest_57; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_58 = digest_58; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_59 = digest_59; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_60 = digest_60; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_61 = digest_61; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_62 = digest_62; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_63 = digest_63; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_64 = digest_64; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_65 = digest_65; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_66 = digest_66; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_67 = digest_67; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_68 = digest_68; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_69 = digest_69; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_70 = digest_70; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_71 = digest_71; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_72 = digest_72; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_73 = digest_73; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_74 = digest_74; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_75 = digest_75; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_76 = digest_76; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_77 = digest_77; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_78 = digest_78; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_arr_79 = digest_79; // @[digest.scala 81:19 315:31]
  assign __m_fill_1_io_off = 32'sh4; // @[digest.scala 81:19 319:31]
  assign __m_fill_1_io_valid = 6'h3f == state ? 1'h0 : _GEN_33710; // @[digest.scala 81:19 63:25]
  assign __m_fill_2_clock = clock;
  assign __m_fill_2_reset = reset;
  assign __m_fill_2_io_value = c; // @[digest.scala 81:19 324:33]
  assign __m_fill_2_io_arr_0 = digest_0; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_1 = digest_1; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_2 = digest_2; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_3 = digest_3; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_4 = digest_4; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_5 = digest_5; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_6 = digest_6; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_7 = digest_7; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_8 = digest_8; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_9 = digest_9; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_10 = digest_10; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_11 = digest_11; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_12 = digest_12; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_13 = digest_13; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_14 = digest_14; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_15 = digest_15; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_16 = digest_16; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_17 = digest_17; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_18 = digest_18; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_19 = digest_19; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_20 = digest_20; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_21 = digest_21; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_22 = digest_22; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_23 = digest_23; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_24 = digest_24; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_25 = digest_25; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_26 = digest_26; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_27 = digest_27; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_28 = digest_28; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_29 = digest_29; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_30 = digest_30; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_31 = digest_31; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_32 = digest_32; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_33 = digest_33; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_34 = digest_34; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_35 = digest_35; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_36 = digest_36; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_37 = digest_37; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_38 = digest_38; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_39 = digest_39; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_40 = digest_40; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_41 = digest_41; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_42 = digest_42; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_43 = digest_43; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_44 = digest_44; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_45 = digest_45; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_46 = digest_46; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_47 = digest_47; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_48 = digest_48; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_49 = digest_49; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_50 = digest_50; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_51 = digest_51; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_52 = digest_52; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_53 = digest_53; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_54 = digest_54; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_55 = digest_55; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_56 = digest_56; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_57 = digest_57; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_58 = digest_58; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_59 = digest_59; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_60 = digest_60; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_61 = digest_61; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_62 = digest_62; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_63 = digest_63; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_64 = digest_64; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_65 = digest_65; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_66 = digest_66; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_67 = digest_67; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_68 = digest_68; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_69 = digest_69; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_70 = digest_70; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_71 = digest_71; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_72 = digest_72; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_73 = digest_73; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_74 = digest_74; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_75 = digest_75; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_76 = digest_76; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_77 = digest_77; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_78 = digest_78; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_arr_79 = digest_79; // @[digest.scala 81:19 325:31]
  assign __m_fill_2_io_off = 32'sh8; // @[digest.scala 81:19 329:31]
  assign __m_fill_2_io_valid = 6'h3f == state ? 1'h0 : _GEN_33793; // @[digest.scala 81:19 68:25]
  assign __m_fill_3_clock = clock;
  assign __m_fill_3_reset = reset;
  assign __m_fill_3_io_value = d; // @[digest.scala 81:19 334:33]
  assign __m_fill_3_io_arr_0 = digest_0; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_1 = digest_1; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_2 = digest_2; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_3 = digest_3; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_4 = digest_4; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_5 = digest_5; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_6 = digest_6; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_7 = digest_7; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_8 = digest_8; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_9 = digest_9; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_10 = digest_10; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_11 = digest_11; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_12 = digest_12; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_13 = digest_13; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_14 = digest_14; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_15 = digest_15; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_16 = digest_16; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_17 = digest_17; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_18 = digest_18; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_19 = digest_19; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_20 = digest_20; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_21 = digest_21; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_22 = digest_22; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_23 = digest_23; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_24 = digest_24; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_25 = digest_25; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_26 = digest_26; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_27 = digest_27; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_28 = digest_28; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_29 = digest_29; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_30 = digest_30; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_31 = digest_31; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_32 = digest_32; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_33 = digest_33; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_34 = digest_34; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_35 = digest_35; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_36 = digest_36; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_37 = digest_37; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_38 = digest_38; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_39 = digest_39; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_40 = digest_40; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_41 = digest_41; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_42 = digest_42; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_43 = digest_43; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_44 = digest_44; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_45 = digest_45; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_46 = digest_46; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_47 = digest_47; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_48 = digest_48; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_49 = digest_49; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_50 = digest_50; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_51 = digest_51; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_52 = digest_52; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_53 = digest_53; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_54 = digest_54; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_55 = digest_55; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_56 = digest_56; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_57 = digest_57; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_58 = digest_58; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_59 = digest_59; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_60 = digest_60; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_61 = digest_61; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_62 = digest_62; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_63 = digest_63; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_64 = digest_64; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_65 = digest_65; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_66 = digest_66; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_67 = digest_67; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_68 = digest_68; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_69 = digest_69; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_70 = digest_70; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_71 = digest_71; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_72 = digest_72; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_73 = digest_73; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_74 = digest_74; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_75 = digest_75; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_76 = digest_76; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_77 = digest_77; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_78 = digest_78; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_arr_79 = digest_79; // @[digest.scala 81:19 335:31]
  assign __m_fill_3_io_off = 32'shc; // @[digest.scala 81:19 339:31]
  assign __m_fill_3_io_valid = 6'h3f == state ? 1'h0 : _GEN_33876; // @[digest.scala 81:19 73:25]
  assign __m_fill_4_clock = clock;
  assign __m_fill_4_reset = reset;
  assign __m_fill_4_io_value = e; // @[digest.scala 81:19 344:33]
  assign __m_fill_4_io_arr_0 = digest_0; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_1 = digest_1; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_2 = digest_2; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_3 = digest_3; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_4 = digest_4; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_5 = digest_5; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_6 = digest_6; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_7 = digest_7; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_8 = digest_8; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_9 = digest_9; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_10 = digest_10; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_11 = digest_11; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_12 = digest_12; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_13 = digest_13; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_14 = digest_14; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_15 = digest_15; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_16 = digest_16; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_17 = digest_17; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_18 = digest_18; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_19 = digest_19; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_20 = digest_20; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_21 = digest_21; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_22 = digest_22; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_23 = digest_23; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_24 = digest_24; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_25 = digest_25; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_26 = digest_26; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_27 = digest_27; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_28 = digest_28; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_29 = digest_29; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_30 = digest_30; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_31 = digest_31; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_32 = digest_32; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_33 = digest_33; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_34 = digest_34; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_35 = digest_35; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_36 = digest_36; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_37 = digest_37; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_38 = digest_38; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_39 = digest_39; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_40 = digest_40; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_41 = digest_41; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_42 = digest_42; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_43 = digest_43; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_44 = digest_44; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_45 = digest_45; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_46 = digest_46; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_47 = digest_47; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_48 = digest_48; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_49 = digest_49; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_50 = digest_50; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_51 = digest_51; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_52 = digest_52; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_53 = digest_53; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_54 = digest_54; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_55 = digest_55; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_56 = digest_56; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_57 = digest_57; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_58 = digest_58; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_59 = digest_59; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_60 = digest_60; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_61 = digest_61; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_62 = digest_62; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_63 = digest_63; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_64 = digest_64; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_65 = digest_65; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_66 = digest_66; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_67 = digest_67; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_68 = digest_68; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_69 = digest_69; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_70 = digest_70; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_71 = digest_71; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_72 = digest_72; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_73 = digest_73; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_74 = digest_74; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_75 = digest_75; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_76 = digest_76; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_77 = digest_77; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_78 = digest_78; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_arr_79 = digest_79; // @[digest.scala 81:19 345:31]
  assign __m_fill_4_io_off = 32'sh10; // @[digest.scala 81:19 349:31]
  assign __m_fill_4_io_valid = 6'h3f == state ? 1'h0 : _GEN_33959; // @[digest.scala 81:19 78:25]
  always @(posedge clock) begin
    if (reset) begin // @[digest.scala 14:24]
      state <= 6'h3f; // @[digest.scala 14:24]
    end else if (6'h3f == state) begin // @[digest.scala 81:19]
      if (io_valid) begin // @[digest.scala 83:25]
        state <= 6'h0;
      end
    end else if (6'h0 == state) begin // @[digest.scala 81:19]
      state <= 6'h1; // @[digest.scala 87:19]
    end else if (6'h1 == state) begin // @[digest.scala 81:19]
      state <= 6'h2; // @[digest.scala 91:19]
    end else begin
      state <= _GEN_31921;
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_0 <= io_bytes_0; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_1 <= io_bytes_1; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_2 <= io_bytes_2; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_3 <= io_bytes_3; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_4 <= io_bytes_4; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_5 <= io_bytes_5; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_6 <= io_bytes_6; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_7 <= io_bytes_7; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_8 <= io_bytes_8; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_9 <= io_bytes_9; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_10 <= io_bytes_10; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_11 <= io_bytes_11; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_12 <= io_bytes_12; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_13 <= io_bytes_13; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_14 <= io_bytes_14; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_15 <= io_bytes_15; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_16 <= io_bytes_16; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_17 <= io_bytes_17; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_18 <= io_bytes_18; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_19 <= io_bytes_19; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_20 <= io_bytes_20; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_21 <= io_bytes_21; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_22 <= io_bytes_22; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_23 <= io_bytes_23; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_24 <= io_bytes_24; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_25 <= io_bytes_25; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_26 <= io_bytes_26; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_27 <= io_bytes_27; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_28 <= io_bytes_28; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_29 <= io_bytes_29; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_30 <= io_bytes_30; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_31 <= io_bytes_31; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_32 <= io_bytes_32; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_33 <= io_bytes_33; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_34 <= io_bytes_34; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_35 <= io_bytes_35; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_36 <= io_bytes_36; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_37 <= io_bytes_37; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_38 <= io_bytes_38; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_39 <= io_bytes_39; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_40 <= io_bytes_40; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_41 <= io_bytes_41; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_42 <= io_bytes_42; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_43 <= io_bytes_43; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_44 <= io_bytes_44; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_45 <= io_bytes_45; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_46 <= io_bytes_46; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_47 <= io_bytes_47; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_48 <= io_bytes_48; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_49 <= io_bytes_49; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_50 <= io_bytes_50; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_51 <= io_bytes_51; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_52 <= io_bytes_52; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_53 <= io_bytes_53; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_54 <= io_bytes_54; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_55 <= io_bytes_55; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_56 <= io_bytes_56; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_57 <= io_bytes_57; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_58 <= io_bytes_58; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_59 <= io_bytes_59; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_60 <= io_bytes_60; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_61 <= io_bytes_61; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_62 <= io_bytes_62; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_63 <= io_bytes_63; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_64 <= io_bytes_64; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_65 <= io_bytes_65; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_66 <= io_bytes_66; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_67 <= io_bytes_67; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_68 <= io_bytes_68; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_69 <= io_bytes_69; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_70 <= io_bytes_70; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_71 <= io_bytes_71; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_72 <= io_bytes_72; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_73 <= io_bytes_73; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_74 <= io_bytes_74; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_75 <= io_bytes_75; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_76 <= io_bytes_76; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_77 <= io_bytes_77; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_78 <= io_bytes_78; // @[digest.scala 20:15]
    end
    if (REG) begin // @[digest.scala 19:29]
      bytes_79 <= io_bytes_79; // @[digest.scala 20:15]
    end
    REG <= ~io_valid; // @[digest.scala 19:18]
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (6'h2 == state) begin // @[digest.scala 81:19]
            i <= 32'sh0; // @[digest.scala 94:15]
          end else begin
            i <= _GEN_31323;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            a <= _GEN_31324;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            b <= _GEN_31325;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            c <= _GEN_31326;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            d <= _GEN_31327;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            e <= _GEN_31328;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            olda <= _GEN_31329;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            oldb <= _GEN_31330;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            oldc <= _GEN_31331;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            oldd <= _GEN_31332;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            olde <= _GEN_31333;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            j <= _GEN_31334;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            t <= _GEN_31418;
          end
        end
      end
    end
    blksLength <= _GEN_33962[31:0];
    temp <= _GEN_33964[31:0];
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_0 <= _GEN_31243;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_1 <= _GEN_31244;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_2 <= _GEN_31245;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_3 <= _GEN_31246;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_4 <= _GEN_31247;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_5 <= _GEN_31248;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_6 <= _GEN_31249;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_7 <= _GEN_31250;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_8 <= _GEN_31251;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_9 <= _GEN_31252;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_10 <= _GEN_31253;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_11 <= _GEN_31254;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_12 <= _GEN_31255;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_13 <= _GEN_31256;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_14 <= _GEN_31257;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_15 <= _GEN_31258;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_16 <= _GEN_31259;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_17 <= _GEN_31260;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_18 <= _GEN_31261;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_19 <= _GEN_31262;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_20 <= _GEN_31263;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_21 <= _GEN_31264;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_22 <= _GEN_31265;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_23 <= _GEN_31266;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_24 <= _GEN_31267;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_25 <= _GEN_31268;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_26 <= _GEN_31269;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_27 <= _GEN_31270;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_28 <= _GEN_31271;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_29 <= _GEN_31272;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_30 <= _GEN_31273;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_31 <= _GEN_31274;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_32 <= _GEN_31275;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_33 <= _GEN_31276;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_34 <= _GEN_31277;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_35 <= _GEN_31278;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_36 <= _GEN_31279;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_37 <= _GEN_31280;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_38 <= _GEN_31281;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_39 <= _GEN_31282;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_40 <= _GEN_31283;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_41 <= _GEN_31284;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_42 <= _GEN_31285;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_43 <= _GEN_31286;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_44 <= _GEN_31287;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_45 <= _GEN_31288;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_46 <= _GEN_31289;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_47 <= _GEN_31290;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_48 <= _GEN_31291;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_49 <= _GEN_31292;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_50 <= _GEN_31293;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_51 <= _GEN_31294;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_52 <= _GEN_31295;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_53 <= _GEN_31296;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_54 <= _GEN_31297;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_55 <= _GEN_31298;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_56 <= _GEN_31299;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_57 <= _GEN_31300;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_58 <= _GEN_31301;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_59 <= _GEN_31302;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_60 <= _GEN_31303;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_61 <= _GEN_31304;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_62 <= _GEN_31305;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_63 <= _GEN_31306;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_64 <= _GEN_31307;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_65 <= _GEN_31308;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_66 <= _GEN_31309;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_67 <= _GEN_31310;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_68 <= _GEN_31311;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_69 <= _GEN_31312;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_70 <= _GEN_31313;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_71 <= _GEN_31314;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_72 <= _GEN_31315;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_73 <= _GEN_31316;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_74 <= _GEN_31317;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_75 <= _GEN_31318;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_76 <= _GEN_31319;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_77 <= _GEN_31320;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_78 <= _GEN_31321;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            blks_79 <= _GEN_31322;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_0 <= _GEN_31335;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_1 <= _GEN_31336;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_2 <= _GEN_31337;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_3 <= _GEN_31338;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_4 <= _GEN_31339;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_5 <= _GEN_31340;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_6 <= _GEN_31341;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_7 <= _GEN_31342;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_8 <= _GEN_31343;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_9 <= _GEN_31344;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_10 <= _GEN_31345;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_11 <= _GEN_31346;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_12 <= _GEN_31347;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_13 <= _GEN_31348;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_14 <= _GEN_31349;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_15 <= _GEN_31350;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_16 <= _GEN_31351;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_17 <= _GEN_31352;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_18 <= _GEN_31353;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_19 <= _GEN_31354;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_20 <= _GEN_31355;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_21 <= _GEN_31356;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_22 <= _GEN_31357;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_23 <= _GEN_31358;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_24 <= _GEN_31359;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_25 <= _GEN_31360;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_26 <= _GEN_31361;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_27 <= _GEN_31362;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_28 <= _GEN_31363;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_29 <= _GEN_31364;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_30 <= _GEN_31365;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_31 <= _GEN_31366;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_32 <= _GEN_31367;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_33 <= _GEN_31368;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_34 <= _GEN_31369;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_35 <= _GEN_31370;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_36 <= _GEN_31371;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_37 <= _GEN_31372;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_38 <= _GEN_31373;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_39 <= _GEN_31374;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_40 <= _GEN_31375;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_41 <= _GEN_31376;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_42 <= _GEN_31377;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_43 <= _GEN_31378;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_44 <= _GEN_31379;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_45 <= _GEN_31380;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_46 <= _GEN_31381;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_47 <= _GEN_31382;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_48 <= _GEN_31383;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_49 <= _GEN_31384;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_50 <= _GEN_31385;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_51 <= _GEN_31386;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_52 <= _GEN_31387;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_53 <= _GEN_31388;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_54 <= _GEN_31389;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_55 <= _GEN_31390;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_56 <= _GEN_31391;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_57 <= _GEN_31392;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_58 <= _GEN_31393;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_59 <= _GEN_31394;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_60 <= _GEN_31395;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_61 <= _GEN_31396;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_62 <= _GEN_31397;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_63 <= _GEN_31398;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_64 <= _GEN_31399;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_65 <= _GEN_31400;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_66 <= _GEN_31401;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_67 <= _GEN_31402;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_68 <= _GEN_31403;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_69 <= _GEN_31404;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_70 <= _GEN_31405;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_71 <= _GEN_31406;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_72 <= _GEN_31407;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_73 <= _GEN_31408;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_74 <= _GEN_31409;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_75 <= _GEN_31410;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_76 <= _GEN_31411;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_77 <= _GEN_31412;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_78 <= _GEN_31413;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            w_79 <= _GEN_31414;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_0 <= _GEN_31506;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_1 <= _GEN_31507;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_2 <= _GEN_31508;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_3 <= _GEN_31509;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_4 <= _GEN_31510;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_5 <= _GEN_31511;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_6 <= _GEN_31512;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_7 <= _GEN_31513;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_8 <= _GEN_31514;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_9 <= _GEN_31515;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_10 <= _GEN_31516;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_11 <= _GEN_31517;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_12 <= _GEN_31518;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_13 <= _GEN_31519;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_14 <= _GEN_31520;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_15 <= _GEN_31521;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_16 <= _GEN_31522;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_17 <= _GEN_31523;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_18 <= _GEN_31524;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_19 <= _GEN_31525;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_20 <= _GEN_31526;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_21 <= _GEN_31527;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_22 <= _GEN_31528;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_23 <= _GEN_31529;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_24 <= _GEN_31530;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_25 <= _GEN_31531;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_26 <= _GEN_31532;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_27 <= _GEN_31533;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_28 <= _GEN_31534;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_29 <= _GEN_31535;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_30 <= _GEN_31536;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_31 <= _GEN_31537;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_32 <= _GEN_31538;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_33 <= _GEN_31539;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_34 <= _GEN_31540;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_35 <= _GEN_31541;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_36 <= _GEN_31542;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_37 <= _GEN_31543;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_38 <= _GEN_31544;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_39 <= _GEN_31545;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_40 <= _GEN_31546;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_41 <= _GEN_31547;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_42 <= _GEN_31548;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_43 <= _GEN_31549;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_44 <= _GEN_31550;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_45 <= _GEN_31551;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_46 <= _GEN_31552;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_47 <= _GEN_31553;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_48 <= _GEN_31554;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_49 <= _GEN_31555;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_50 <= _GEN_31556;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_51 <= _GEN_31557;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_52 <= _GEN_31558;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_53 <= _GEN_31559;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_54 <= _GEN_31560;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_55 <= _GEN_31561;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_56 <= _GEN_31562;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_57 <= _GEN_31563;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_58 <= _GEN_31564;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_59 <= _GEN_31565;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_60 <= _GEN_31566;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_61 <= _GEN_31567;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_62 <= _GEN_31568;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_63 <= _GEN_31569;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_64 <= _GEN_31570;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_65 <= _GEN_31571;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_66 <= _GEN_31572;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_67 <= _GEN_31573;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_68 <= _GEN_31574;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_69 <= _GEN_31575;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_70 <= _GEN_31576;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_71 <= _GEN_31577;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_72 <= _GEN_31578;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_73 <= _GEN_31579;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_74 <= _GEN_31580;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_75 <= _GEN_31581;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_76 <= _GEN_31582;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_77 <= _GEN_31583;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_78 <= _GEN_31584;
          end
        end
      end
    end
    if (!(6'h3f == state)) begin // @[digest.scala 81:19]
      if (!(6'h0 == state)) begin // @[digest.scala 81:19]
        if (!(6'h1 == state)) begin // @[digest.scala 81:19]
          if (!(6'h2 == state)) begin // @[digest.scala 81:19]
            digest_79 <= _GEN_31585;
          end
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  bytes_0 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  bytes_1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  bytes_2 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  bytes_3 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  bytes_4 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  bytes_5 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  bytes_6 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  bytes_7 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  bytes_8 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  bytes_9 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  bytes_10 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  bytes_11 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  bytes_12 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  bytes_13 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  bytes_14 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  bytes_15 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  bytes_16 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  bytes_17 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  bytes_18 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  bytes_19 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  bytes_20 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  bytes_21 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  bytes_22 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  bytes_23 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  bytes_24 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  bytes_25 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  bytes_26 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  bytes_27 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  bytes_28 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  bytes_29 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  bytes_30 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  bytes_31 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  bytes_32 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  bytes_33 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  bytes_34 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  bytes_35 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  bytes_36 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  bytes_37 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  bytes_38 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  bytes_39 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  bytes_40 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  bytes_41 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  bytes_42 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  bytes_43 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  bytes_44 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  bytes_45 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  bytes_46 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  bytes_47 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  bytes_48 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  bytes_49 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  bytes_50 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  bytes_51 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  bytes_52 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  bytes_53 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  bytes_54 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  bytes_55 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  bytes_56 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  bytes_57 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  bytes_58 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  bytes_59 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  bytes_60 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  bytes_61 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  bytes_62 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  bytes_63 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  bytes_64 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  bytes_65 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  bytes_66 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  bytes_67 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  bytes_68 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  bytes_69 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  bytes_70 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  bytes_71 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  bytes_72 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  bytes_73 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  bytes_74 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  bytes_75 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  bytes_76 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  bytes_77 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  bytes_78 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  bytes_79 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  REG = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  i = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  a = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  b = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  c = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  d = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  e = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  olda = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  oldb = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  oldc = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  oldd = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  olde = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  j = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  t = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  blksLength = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  temp = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  blks_0 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  blks_1 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  blks_2 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  blks_3 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  blks_4 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  blks_5 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  blks_6 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  blks_7 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  blks_8 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  blks_9 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  blks_10 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  blks_11 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  blks_12 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  blks_13 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  blks_14 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  blks_15 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  blks_16 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  blks_17 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  blks_18 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  blks_19 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  blks_20 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  blks_21 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  blks_22 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  blks_23 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  blks_24 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  blks_25 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  blks_26 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  blks_27 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  blks_28 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  blks_29 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  blks_30 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  blks_31 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  blks_32 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  blks_33 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  blks_34 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  blks_35 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  blks_36 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  blks_37 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  blks_38 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  blks_39 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  blks_40 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  blks_41 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  blks_42 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  blks_43 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  blks_44 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  blks_45 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  blks_46 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  blks_47 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  blks_48 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  blks_49 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  blks_50 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  blks_51 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  blks_52 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  blks_53 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  blks_54 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  blks_55 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  blks_56 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  blks_57 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  blks_58 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  blks_59 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  blks_60 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  blks_61 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  blks_62 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  blks_63 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  blks_64 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  blks_65 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  blks_66 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  blks_67 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  blks_68 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  blks_69 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  blks_70 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  blks_71 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  blks_72 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  blks_73 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  blks_74 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  blks_75 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  blks_76 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  blks_77 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  blks_78 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  blks_79 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  w_0 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  w_1 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  w_2 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  w_3 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  w_4 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  w_5 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  w_6 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  w_7 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  w_8 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  w_9 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  w_10 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  w_11 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  w_12 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  w_13 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  w_14 = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  w_15 = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  w_16 = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  w_17 = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  w_18 = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  w_19 = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  w_20 = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  w_21 = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  w_22 = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  w_23 = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  w_24 = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  w_25 = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  w_26 = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  w_27 = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  w_28 = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  w_29 = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  w_30 = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  w_31 = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  w_32 = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  w_33 = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  w_34 = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  w_35 = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  w_36 = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  w_37 = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  w_38 = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  w_39 = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  w_40 = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  w_41 = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  w_42 = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  w_43 = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  w_44 = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  w_45 = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  w_46 = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  w_47 = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  w_48 = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  w_49 = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  w_50 = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  w_51 = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  w_52 = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  w_53 = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  w_54 = _RAND_231[31:0];
  _RAND_232 = {1{`RANDOM}};
  w_55 = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  w_56 = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  w_57 = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  w_58 = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  w_59 = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  w_60 = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  w_61 = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  w_62 = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  w_63 = _RAND_240[31:0];
  _RAND_241 = {1{`RANDOM}};
  w_64 = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  w_65 = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  w_66 = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  w_67 = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  w_68 = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  w_69 = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  w_70 = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  w_71 = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  w_72 = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  w_73 = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  w_74 = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  w_75 = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  w_76 = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  w_77 = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  w_78 = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  w_79 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  digest_0 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  digest_1 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  digest_2 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  digest_3 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  digest_4 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  digest_5 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  digest_6 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  digest_7 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  digest_8 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  digest_9 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  digest_10 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  digest_11 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  digest_12 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  digest_13 = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  digest_14 = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  digest_15 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  digest_16 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  digest_17 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  digest_18 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  digest_19 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  digest_20 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  digest_21 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  digest_22 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  digest_23 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  digest_24 = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  digest_25 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  digest_26 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  digest_27 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  digest_28 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  digest_29 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  digest_30 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  digest_31 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  digest_32 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  digest_33 = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  digest_34 = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  digest_35 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  digest_36 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  digest_37 = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  digest_38 = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  digest_39 = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  digest_40 = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  digest_41 = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  digest_42 = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  digest_43 = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  digest_44 = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  digest_45 = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  digest_46 = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  digest_47 = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  digest_48 = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  digest_49 = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  digest_50 = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  digest_51 = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  digest_52 = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  digest_53 = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  digest_54 = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  digest_55 = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  digest_56 = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  digest_57 = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  digest_58 = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  digest_59 = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  digest_60 = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  digest_61 = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  digest_62 = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  digest_63 = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  digest_64 = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  digest_65 = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  digest_66 = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  digest_67 = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  digest_68 = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  digest_69 = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  digest_70 = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  digest_71 = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  digest_72 = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  digest_73 = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  digest_74 = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  digest_75 = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  digest_76 = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  digest_77 = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  digest_78 = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  digest_79 = _RAND_336[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule