[info] welcome to sbt 1.9.7 (Ubuntu Java 11.0.19)
[info] loading settings for project chisel-template-build from plugins.sbt ...
[info] loading project definition from /share/git_dir/chisel-template/project
[info] loading settings for project chisel-template from build.sbt ...
[info] set current project to chisel-template (in build file:/share/git_dir/chisel-template/)
[warn] sbt 0.13 shell syntax is deprecated; use slash syntax instead: Test / runMain
[info] compiling 1 Scala source to /share/git_dir/chisel-template/target/scala-2.12/test-classes ...
[info] done compiling
[warn] multiple main classes detected: run 'show discoveredMainClasses' to see the list
[info] running AXIWrapperChisel.AXIWrapperChiselInsertSortVerilogGeneration 
module insertSort(
  input         clock,
  input         reset,
  input  [31:0] io_array_0,
  input  [31:0] io_array_1,
  input  [31:0] io_array_2,
  input  [31:0] io_array_3,
  input  [31:0] io_array_4,
  input  [31:0] io_array_5,
  input  [31:0] io_array_6,
  input  [31:0] io_array_7,
  input  [31:0] io_array_8,
  input  [31:0] io_array_9,
  input  [31:0] io_array_10,
  input  [31:0] io_array_11,
  input  [31:0] io_array_12,
  input  [31:0] io_array_13,
  input  [31:0] io_array_14,
  input  [31:0] io_array_15,
  input  [31:0] io_array_16,
  input  [31:0] io_array_17,
  input  [31:0] io_array_18,
  input  [31:0] io_array_19,
  input         io_valid,
  output [31:0] io_array_out_0,
  output [31:0] io_array_out_1,
  output [31:0] io_array_out_2,
  output [31:0] io_array_out_3,
  output [31:0] io_array_out_4,
  output [31:0] io_array_out_5,
  output [31:0] io_array_out_6,
  output [31:0] io_array_out_7,
  output [31:0] io_array_out_8,
  output [31:0] io_array_out_9,
  output [31:0] io_array_out_10,
  output [31:0] io_array_out_11,
  output [31:0] io_array_out_12,
  output [31:0] io_array_out_13,
  output [31:0] io_array_out_14,
  output [31:0] io_array_out_15,
  output [31:0] io_array_out_16,
  output [31:0] io_array_out_17,
  output [31:0] io_array_out_18,
  output [31:0] io_array_out_19,
  output        io_ready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] state; // @[insertSort.scala 13:24]
  wire [3:0] _GEN_0 = reset ? 4'hf : state; // @[insertSort.scala 14:26 15:15 13:24]
  reg [31:0] array_0; // @[insertSort.scala 17:20]
  reg [31:0] array_1; // @[insertSort.scala 17:20]
  reg [31:0] array_2; // @[insertSort.scala 17:20]
  reg [31:0] array_3; // @[insertSort.scala 17:20]
  reg [31:0] array_4; // @[insertSort.scala 17:20]
  reg [31:0] array_5; // @[insertSort.scala 17:20]
  reg [31:0] array_6; // @[insertSort.scala 17:20]
  reg [31:0] array_7; // @[insertSort.scala 17:20]
  reg [31:0] array_8; // @[insertSort.scala 17:20]
  reg [31:0] array_9; // @[insertSort.scala 17:20]
  reg [31:0] array_10; // @[insertSort.scala 17:20]
  reg [31:0] array_11; // @[insertSort.scala 17:20]
  reg [31:0] array_12; // @[insertSort.scala 17:20]
  reg [31:0] array_13; // @[insertSort.scala 17:20]
  reg [31:0] array_14; // @[insertSort.scala 17:20]
  reg [31:0] array_15; // @[insertSort.scala 17:20]
  reg [31:0] array_16; // @[insertSort.scala 17:20]
  reg [31:0] array_17; // @[insertSort.scala 17:20]
  reg [31:0] array_18; // @[insertSort.scala 17:20]
  reg [31:0] array_19; // @[insertSort.scala 17:20]
  reg [31:0] array_20; // @[insertSort.scala 17:20]
  reg [31:0] array_21; // @[insertSort.scala 17:20]
  reg [31:0] array_22; // @[insertSort.scala 17:20]
  reg [31:0] array_23; // @[insertSort.scala 17:20]
  reg [31:0] array_24; // @[insertSort.scala 17:20]
  reg [31:0] array_25; // @[insertSort.scala 17:20]
  reg [31:0] array_26; // @[insertSort.scala 17:20]
  reg [31:0] array_27; // @[insertSort.scala 17:20]
  reg [31:0] array_28; // @[insertSort.scala 17:20]
  reg [31:0] array_29; // @[insertSort.scala 17:20]
  reg [31:0] array_30; // @[insertSort.scala 17:20]
  reg [31:0] array_31; // @[insertSort.scala 17:20]
  reg [31:0] array_32; // @[insertSort.scala 17:20]
  reg [31:0] array_33; // @[insertSort.scala 17:20]
  reg [31:0] array_34; // @[insertSort.scala 17:20]
  reg [31:0] array_35; // @[insertSort.scala 17:20]
  reg [31:0] array_36; // @[insertSort.scala 17:20]
  reg [31:0] array_37; // @[insertSort.scala 17:20]
  reg [31:0] array_38; // @[insertSort.scala 17:20]
  reg [31:0] array_39; // @[insertSort.scala 17:20]
  reg [31:0] array_40; // @[insertSort.scala 17:20]
  reg [31:0] array_41; // @[insertSort.scala 17:20]
  reg [31:0] array_42; // @[insertSort.scala 17:20]
  reg [31:0] array_43; // @[insertSort.scala 17:20]
  reg [31:0] array_44; // @[insertSort.scala 17:20]
  reg [31:0] array_45; // @[insertSort.scala 17:20]
  reg [31:0] array_46; // @[insertSort.scala 17:20]
  reg [31:0] array_47; // @[insertSort.scala 17:20]
  reg [31:0] array_48; // @[insertSort.scala 17:20]
  reg [31:0] array_49; // @[insertSort.scala 17:20]
  reg [31:0] array_50; // @[insertSort.scala 17:20]
  reg [31:0] array_51; // @[insertSort.scala 17:20]
  reg [31:0] array_52; // @[insertSort.scala 17:20]
  reg [31:0] array_53; // @[insertSort.scala 17:20]
  reg [31:0] array_54; // @[insertSort.scala 17:20]
  reg [31:0] array_55; // @[insertSort.scala 17:20]
  reg [31:0] array_56; // @[insertSort.scala 17:20]
  reg [31:0] array_57; // @[insertSort.scala 17:20]
  reg [31:0] array_58; // @[insertSort.scala 17:20]
  reg [31:0] array_59; // @[insertSort.scala 17:20]
  reg [31:0] array_60; // @[insertSort.scala 17:20]
  reg [31:0] array_61; // @[insertSort.scala 17:20]
  reg [31:0] array_62; // @[insertSort.scala 17:20]
  reg [31:0] array_63; // @[insertSort.scala 17:20]
  reg [31:0] array_64; // @[insertSort.scala 17:20]
  reg [31:0] array_65; // @[insertSort.scala 17:20]
  reg [31:0] array_66; // @[insertSort.scala 17:20]
  reg [31:0] array_67; // @[insertSort.scala 17:20]
  reg [31:0] array_68; // @[insertSort.scala 17:20]
  reg [31:0] array_69; // @[insertSort.scala 17:20]
  reg [31:0] array_70; // @[insertSort.scala 17:20]
  reg [31:0] array_71; // @[insertSort.scala 17:20]
  reg [31:0] array_72; // @[insertSort.scala 17:20]
  reg [31:0] array_73; // @[insertSort.scala 17:20]
  reg [31:0] array_74; // @[insertSort.scala 17:20]
  reg [31:0] array_75; // @[insertSort.scala 17:20]
  reg [31:0] array_76; // @[insertSort.scala 17:20]
  reg [31:0] array_77; // @[insertSort.scala 17:20]
  reg [31:0] array_78; // @[insertSort.scala 17:20]
  reg [31:0] array_79; // @[insertSort.scala 17:20]
  reg  REG; // @[insertSort.scala 18:17]
  wire [31:0] _GEN_1 = REG ? $signed(io_array_0) : $signed(array_0); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_2 = REG ? $signed(io_array_1) : $signed(array_1); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_3 = REG ? $signed(io_array_2) : $signed(array_2); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_4 = REG ? $signed(io_array_3) : $signed(array_3); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_5 = REG ? $signed(io_array_4) : $signed(array_4); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_6 = REG ? $signed(io_array_5) : $signed(array_5); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_7 = REG ? $signed(io_array_6) : $signed(array_6); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_8 = REG ? $signed(io_array_7) : $signed(array_7); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_9 = REG ? $signed(io_array_8) : $signed(array_8); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_10 = REG ? $signed(io_array_9) : $signed(array_9); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_11 = REG ? $signed(io_array_10) : $signed(array_10); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_12 = REG ? $signed(io_array_11) : $signed(array_11); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_13 = REG ? $signed(io_array_12) : $signed(array_12); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_14 = REG ? $signed(io_array_13) : $signed(array_13); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_15 = REG ? $signed(io_array_14) : $signed(array_14); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_16 = REG ? $signed(io_array_15) : $signed(array_15); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_17 = REG ? $signed(io_array_16) : $signed(array_16); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_18 = REG ? $signed(io_array_17) : $signed(array_17); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_19 = REG ? $signed(io_array_18) : $signed(array_18); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_20 = REG ? $signed(io_array_19) : $signed(array_19); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_21 = REG ? $signed(32'sh0) : $signed(array_20); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_22 = REG ? $signed(32'sh0) : $signed(array_21); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_23 = REG ? $signed(32'sh0) : $signed(array_22); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_24 = REG ? $signed(32'sh0) : $signed(array_23); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_25 = REG ? $signed(32'sh0) : $signed(array_24); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_26 = REG ? $signed(32'sh0) : $signed(array_25); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_27 = REG ? $signed(32'sh0) : $signed(array_26); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_28 = REG ? $signed(32'sh0) : $signed(array_27); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_29 = REG ? $signed(32'sh0) : $signed(array_28); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_30 = REG ? $signed(32'sh0) : $signed(array_29); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_31 = REG ? $signed(32'sh0) : $signed(array_30); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_32 = REG ? $signed(32'sh0) : $signed(array_31); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_33 = REG ? $signed(32'sh0) : $signed(array_32); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_34 = REG ? $signed(32'sh0) : $signed(array_33); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_35 = REG ? $signed(32'sh0) : $signed(array_34); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_36 = REG ? $signed(32'sh0) : $signed(array_35); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_37 = REG ? $signed(32'sh0) : $signed(array_36); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_38 = REG ? $signed(32'sh0) : $signed(array_37); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_39 = REG ? $signed(32'sh0) : $signed(array_38); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_40 = REG ? $signed(32'sh0) : $signed(array_39); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_41 = REG ? $signed(32'sh0) : $signed(array_40); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_42 = REG ? $signed(32'sh0) : $signed(array_41); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_43 = REG ? $signed(32'sh0) : $signed(array_42); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_44 = REG ? $signed(32'sh0) : $signed(array_43); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_45 = REG ? $signed(32'sh0) : $signed(array_44); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_46 = REG ? $signed(32'sh0) : $signed(array_45); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_47 = REG ? $signed(32'sh0) : $signed(array_46); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_48 = REG ? $signed(32'sh0) : $signed(array_47); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_49 = REG ? $signed(32'sh0) : $signed(array_48); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_50 = REG ? $signed(32'sh0) : $signed(array_49); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_51 = REG ? $signed(32'sh0) : $signed(array_50); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_52 = REG ? $signed(32'sh0) : $signed(array_51); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_53 = REG ? $signed(32'sh0) : $signed(array_52); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_54 = REG ? $signed(32'sh0) : $signed(array_53); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_55 = REG ? $signed(32'sh0) : $signed(array_54); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_56 = REG ? $signed(32'sh0) : $signed(array_55); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_57 = REG ? $signed(32'sh0) : $signed(array_56); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_58 = REG ? $signed(32'sh0) : $signed(array_57); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_59 = REG ? $signed(32'sh0) : $signed(array_58); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_60 = REG ? $signed(32'sh0) : $signed(array_59); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_61 = REG ? $signed(32'sh0) : $signed(array_60); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_62 = REG ? $signed(32'sh0) : $signed(array_61); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_63 = REG ? $signed(32'sh0) : $signed(array_62); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_64 = REG ? $signed(32'sh0) : $signed(array_63); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_65 = REG ? $signed(32'sh0) : $signed(array_64); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_66 = REG ? $signed(32'sh0) : $signed(array_65); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_67 = REG ? $signed(32'sh0) : $signed(array_66); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_68 = REG ? $signed(32'sh0) : $signed(array_67); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_69 = REG ? $signed(32'sh0) : $signed(array_68); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_70 = REG ? $signed(32'sh0) : $signed(array_69); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_71 = REG ? $signed(32'sh0) : $signed(array_70); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_72 = REG ? $signed(32'sh0) : $signed(array_71); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_73 = REG ? $signed(32'sh0) : $signed(array_72); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_74 = REG ? $signed(32'sh0) : $signed(array_73); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_75 = REG ? $signed(32'sh0) : $signed(array_74); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_76 = REG ? $signed(32'sh0) : $signed(array_75); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_77 = REG ? $signed(32'sh0) : $signed(array_76); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_78 = REG ? $signed(32'sh0) : $signed(array_77); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_79 = REG ? $signed(32'sh0) : $signed(array_78); // @[insertSort.scala 18:29 19:15 17:20]
  wire [31:0] _GEN_80 = REG ? $signed(32'sh0) : $signed(array_79); // @[insertSort.scala 18:29 19:15 17:20]
  reg [31:0] i; // @[insertSort.scala 22:16]
  reg [31:0] key; // @[insertSort.scala 23:18]
  reg [31:0] j; // @[insertSort.scala 24:16]
  wire [3:0] _state_T_2 = $signed(i) < 32'sha ? 4'h2 : 4'hc; // @[insertSort.scala 35:25]
  wire [31:0] _key_T = i; // @[insertSort.scala 38:36]
  wire [31:0] _GEN_82 = 7'h1 == _key_T[6:0] ? $signed(array_1) : $signed(array_0); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_83 = 7'h2 == _key_T[6:0] ? $signed(array_2) : $signed(_GEN_82); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_84 = 7'h3 == _key_T[6:0] ? $signed(array_3) : $signed(_GEN_83); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_85 = 7'h4 == _key_T[6:0] ? $signed(array_4) : $signed(_GEN_84); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_86 = 7'h5 == _key_T[6:0] ? $signed(array_5) : $signed(_GEN_85); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_87 = 7'h6 == _key_T[6:0] ? $signed(array_6) : $signed(_GEN_86); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_88 = 7'h7 == _key_T[6:0] ? $signed(array_7) : $signed(_GEN_87); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_89 = 7'h8 == _key_T[6:0] ? $signed(array_8) : $signed(_GEN_88); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_90 = 7'h9 == _key_T[6:0] ? $signed(array_9) : $signed(_GEN_89); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_91 = 7'ha == _key_T[6:0] ? $signed(array_10) : $signed(_GEN_90); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_92 = 7'hb == _key_T[6:0] ? $signed(array_11) : $signed(_GEN_91); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_93 = 7'hc == _key_T[6:0] ? $signed(array_12) : $signed(_GEN_92); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_94 = 7'hd == _key_T[6:0] ? $signed(array_13) : $signed(_GEN_93); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_95 = 7'he == _key_T[6:0] ? $signed(array_14) : $signed(_GEN_94); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_96 = 7'hf == _key_T[6:0] ? $signed(array_15) : $signed(_GEN_95); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_97 = 7'h10 == _key_T[6:0] ? $signed(array_16) : $signed(_GEN_96); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_98 = 7'h11 == _key_T[6:0] ? $signed(array_17) : $signed(_GEN_97); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_99 = 7'h12 == _key_T[6:0] ? $signed(array_18) : $signed(_GEN_98); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_100 = 7'h13 == _key_T[6:0] ? $signed(array_19) : $signed(_GEN_99); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_101 = 7'h14 == _key_T[6:0] ? $signed(array_20) : $signed(_GEN_100); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_102 = 7'h15 == _key_T[6:0] ? $signed(array_21) : $signed(_GEN_101); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_103 = 7'h16 == _key_T[6:0] ? $signed(array_22) : $signed(_GEN_102); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_104 = 7'h17 == _key_T[6:0] ? $signed(array_23) : $signed(_GEN_103); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_105 = 7'h18 == _key_T[6:0] ? $signed(array_24) : $signed(_GEN_104); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_106 = 7'h19 == _key_T[6:0] ? $signed(array_25) : $signed(_GEN_105); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_107 = 7'h1a == _key_T[6:0] ? $signed(array_26) : $signed(_GEN_106); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_108 = 7'h1b == _key_T[6:0] ? $signed(array_27) : $signed(_GEN_107); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_109 = 7'h1c == _key_T[6:0] ? $signed(array_28) : $signed(_GEN_108); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_110 = 7'h1d == _key_T[6:0] ? $signed(array_29) : $signed(_GEN_109); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_111 = 7'h1e == _key_T[6:0] ? $signed(array_30) : $signed(_GEN_110); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_112 = 7'h1f == _key_T[6:0] ? $signed(array_31) : $signed(_GEN_111); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_113 = 7'h20 == _key_T[6:0] ? $signed(array_32) : $signed(_GEN_112); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_114 = 7'h21 == _key_T[6:0] ? $signed(array_33) : $signed(_GEN_113); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_115 = 7'h22 == _key_T[6:0] ? $signed(array_34) : $signed(_GEN_114); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_116 = 7'h23 == _key_T[6:0] ? $signed(array_35) : $signed(_GEN_115); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_117 = 7'h24 == _key_T[6:0] ? $signed(array_36) : $signed(_GEN_116); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_118 = 7'h25 == _key_T[6:0] ? $signed(array_37) : $signed(_GEN_117); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_119 = 7'h26 == _key_T[6:0] ? $signed(array_38) : $signed(_GEN_118); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_120 = 7'h27 == _key_T[6:0] ? $signed(array_39) : $signed(_GEN_119); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_121 = 7'h28 == _key_T[6:0] ? $signed(array_40) : $signed(_GEN_120); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_122 = 7'h29 == _key_T[6:0] ? $signed(array_41) : $signed(_GEN_121); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_123 = 7'h2a == _key_T[6:0] ? $signed(array_42) : $signed(_GEN_122); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_124 = 7'h2b == _key_T[6:0] ? $signed(array_43) : $signed(_GEN_123); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_125 = 7'h2c == _key_T[6:0] ? $signed(array_44) : $signed(_GEN_124); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_126 = 7'h2d == _key_T[6:0] ? $signed(array_45) : $signed(_GEN_125); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_127 = 7'h2e == _key_T[6:0] ? $signed(array_46) : $signed(_GEN_126); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_128 = 7'h2f == _key_T[6:0] ? $signed(array_47) : $signed(_GEN_127); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_129 = 7'h30 == _key_T[6:0] ? $signed(array_48) : $signed(_GEN_128); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_130 = 7'h31 == _key_T[6:0] ? $signed(array_49) : $signed(_GEN_129); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_131 = 7'h32 == _key_T[6:0] ? $signed(array_50) : $signed(_GEN_130); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_132 = 7'h33 == _key_T[6:0] ? $signed(array_51) : $signed(_GEN_131); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_133 = 7'h34 == _key_T[6:0] ? $signed(array_52) : $signed(_GEN_132); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_134 = 7'h35 == _key_T[6:0] ? $signed(array_53) : $signed(_GEN_133); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_135 = 7'h36 == _key_T[6:0] ? $signed(array_54) : $signed(_GEN_134); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_136 = 7'h37 == _key_T[6:0] ? $signed(array_55) : $signed(_GEN_135); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_137 = 7'h38 == _key_T[6:0] ? $signed(array_56) : $signed(_GEN_136); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_138 = 7'h39 == _key_T[6:0] ? $signed(array_57) : $signed(_GEN_137); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_139 = 7'h3a == _key_T[6:0] ? $signed(array_58) : $signed(_GEN_138); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_140 = 7'h3b == _key_T[6:0] ? $signed(array_59) : $signed(_GEN_139); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_141 = 7'h3c == _key_T[6:0] ? $signed(array_60) : $signed(_GEN_140); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_142 = 7'h3d == _key_T[6:0] ? $signed(array_61) : $signed(_GEN_141); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_143 = 7'h3e == _key_T[6:0] ? $signed(array_62) : $signed(_GEN_142); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_144 = 7'h3f == _key_T[6:0] ? $signed(array_63) : $signed(_GEN_143); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_145 = 7'h40 == _key_T[6:0] ? $signed(array_64) : $signed(_GEN_144); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_146 = 7'h41 == _key_T[6:0] ? $signed(array_65) : $signed(_GEN_145); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_147 = 7'h42 == _key_T[6:0] ? $signed(array_66) : $signed(_GEN_146); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_148 = 7'h43 == _key_T[6:0] ? $signed(array_67) : $signed(_GEN_147); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_149 = 7'h44 == _key_T[6:0] ? $signed(array_68) : $signed(_GEN_148); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_150 = 7'h45 == _key_T[6:0] ? $signed(array_69) : $signed(_GEN_149); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_151 = 7'h46 == _key_T[6:0] ? $signed(array_70) : $signed(_GEN_150); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_152 = 7'h47 == _key_T[6:0] ? $signed(array_71) : $signed(_GEN_151); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_153 = 7'h48 == _key_T[6:0] ? $signed(array_72) : $signed(_GEN_152); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_154 = 7'h49 == _key_T[6:0] ? $signed(array_73) : $signed(_GEN_153); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_155 = 7'h4a == _key_T[6:0] ? $signed(array_74) : $signed(_GEN_154); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_156 = 7'h4b == _key_T[6:0] ? $signed(array_75) : $signed(_GEN_155); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_157 = 7'h4c == _key_T[6:0] ? $signed(array_76) : $signed(_GEN_156); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_158 = 7'h4d == _key_T[6:0] ? $signed(array_77) : $signed(_GEN_157); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_159 = 7'h4e == _key_T[6:0] ? $signed(array_78) : $signed(_GEN_158); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _GEN_160 = 7'h4f == _key_T[6:0] ? $signed(array_79) : $signed(_GEN_159); // @[insertSort.scala 38:{17,17}]
  wire [31:0] _j_T_2 = $signed(i) - 32'sh1; // @[insertSort.scala 42:20]
  wire [31:0] _state_T_4 = j; // @[insertSort.scala 46:60]
  wire [31:0] _GEN_162 = 7'h1 == _state_T_4[6:0] ? $signed(array_1) : $signed(array_0); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_163 = 7'h2 == _state_T_4[6:0] ? $signed(array_2) : $signed(_GEN_162); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_164 = 7'h3 == _state_T_4[6:0] ? $signed(array_3) : $signed(_GEN_163); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_165 = 7'h4 == _state_T_4[6:0] ? $signed(array_4) : $signed(_GEN_164); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_166 = 7'h5 == _state_T_4[6:0] ? $signed(array_5) : $signed(_GEN_165); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_167 = 7'h6 == _state_T_4[6:0] ? $signed(array_6) : $signed(_GEN_166); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_168 = 7'h7 == _state_T_4[6:0] ? $signed(array_7) : $signed(_GEN_167); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_169 = 7'h8 == _state_T_4[6:0] ? $signed(array_8) : $signed(_GEN_168); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_170 = 7'h9 == _state_T_4[6:0] ? $signed(array_9) : $signed(_GEN_169); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_171 = 7'ha == _state_T_4[6:0] ? $signed(array_10) : $signed(_GEN_170); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_172 = 7'hb == _state_T_4[6:0] ? $signed(array_11) : $signed(_GEN_171); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_173 = 7'hc == _state_T_4[6:0] ? $signed(array_12) : $signed(_GEN_172); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_174 = 7'hd == _state_T_4[6:0] ? $signed(array_13) : $signed(_GEN_173); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_175 = 7'he == _state_T_4[6:0] ? $signed(array_14) : $signed(_GEN_174); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_176 = 7'hf == _state_T_4[6:0] ? $signed(array_15) : $signed(_GEN_175); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_177 = 7'h10 == _state_T_4[6:0] ? $signed(array_16) : $signed(_GEN_176); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_178 = 7'h11 == _state_T_4[6:0] ? $signed(array_17) : $signed(_GEN_177); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_179 = 7'h12 == _state_T_4[6:0] ? $signed(array_18) : $signed(_GEN_178); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_180 = 7'h13 == _state_T_4[6:0] ? $signed(array_19) : $signed(_GEN_179); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_181 = 7'h14 == _state_T_4[6:0] ? $signed(array_20) : $signed(_GEN_180); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_182 = 7'h15 == _state_T_4[6:0] ? $signed(array_21) : $signed(_GEN_181); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_183 = 7'h16 == _state_T_4[6:0] ? $signed(array_22) : $signed(_GEN_182); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_184 = 7'h17 == _state_T_4[6:0] ? $signed(array_23) : $signed(_GEN_183); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_185 = 7'h18 == _state_T_4[6:0] ? $signed(array_24) : $signed(_GEN_184); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_186 = 7'h19 == _state_T_4[6:0] ? $signed(array_25) : $signed(_GEN_185); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_187 = 7'h1a == _state_T_4[6:0] ? $signed(array_26) : $signed(_GEN_186); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_188 = 7'h1b == _state_T_4[6:0] ? $signed(array_27) : $signed(_GEN_187); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_189 = 7'h1c == _state_T_4[6:0] ? $signed(array_28) : $signed(_GEN_188); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_190 = 7'h1d == _state_T_4[6:0] ? $signed(array_29) : $signed(_GEN_189); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_191 = 7'h1e == _state_T_4[6:0] ? $signed(array_30) : $signed(_GEN_190); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_192 = 7'h1f == _state_T_4[6:0] ? $signed(array_31) : $signed(_GEN_191); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_193 = 7'h20 == _state_T_4[6:0] ? $signed(array_32) : $signed(_GEN_192); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_194 = 7'h21 == _state_T_4[6:0] ? $signed(array_33) : $signed(_GEN_193); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_195 = 7'h22 == _state_T_4[6:0] ? $signed(array_34) : $signed(_GEN_194); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_196 = 7'h23 == _state_T_4[6:0] ? $signed(array_35) : $signed(_GEN_195); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_197 = 7'h24 == _state_T_4[6:0] ? $signed(array_36) : $signed(_GEN_196); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_198 = 7'h25 == _state_T_4[6:0] ? $signed(array_37) : $signed(_GEN_197); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_199 = 7'h26 == _state_T_4[6:0] ? $signed(array_38) : $signed(_GEN_198); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_200 = 7'h27 == _state_T_4[6:0] ? $signed(array_39) : $signed(_GEN_199); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_201 = 7'h28 == _state_T_4[6:0] ? $signed(array_40) : $signed(_GEN_200); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_202 = 7'h29 == _state_T_4[6:0] ? $signed(array_41) : $signed(_GEN_201); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_203 = 7'h2a == _state_T_4[6:0] ? $signed(array_42) : $signed(_GEN_202); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_204 = 7'h2b == _state_T_4[6:0] ? $signed(array_43) : $signed(_GEN_203); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_205 = 7'h2c == _state_T_4[6:0] ? $signed(array_44) : $signed(_GEN_204); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_206 = 7'h2d == _state_T_4[6:0] ? $signed(array_45) : $signed(_GEN_205); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_207 = 7'h2e == _state_T_4[6:0] ? $signed(array_46) : $signed(_GEN_206); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_208 = 7'h2f == _state_T_4[6:0] ? $signed(array_47) : $signed(_GEN_207); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_209 = 7'h30 == _state_T_4[6:0] ? $signed(array_48) : $signed(_GEN_208); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_210 = 7'h31 == _state_T_4[6:0] ? $signed(array_49) : $signed(_GEN_209); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_211 = 7'h32 == _state_T_4[6:0] ? $signed(array_50) : $signed(_GEN_210); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_212 = 7'h33 == _state_T_4[6:0] ? $signed(array_51) : $signed(_GEN_211); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_213 = 7'h34 == _state_T_4[6:0] ? $signed(array_52) : $signed(_GEN_212); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_214 = 7'h35 == _state_T_4[6:0] ? $signed(array_53) : $signed(_GEN_213); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_215 = 7'h36 == _state_T_4[6:0] ? $signed(array_54) : $signed(_GEN_214); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_216 = 7'h37 == _state_T_4[6:0] ? $signed(array_55) : $signed(_GEN_215); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_217 = 7'h38 == _state_T_4[6:0] ? $signed(array_56) : $signed(_GEN_216); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_218 = 7'h39 == _state_T_4[6:0] ? $signed(array_57) : $signed(_GEN_217); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_219 = 7'h3a == _state_T_4[6:0] ? $signed(array_58) : $signed(_GEN_218); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_220 = 7'h3b == _state_T_4[6:0] ? $signed(array_59) : $signed(_GEN_219); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_221 = 7'h3c == _state_T_4[6:0] ? $signed(array_60) : $signed(_GEN_220); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_222 = 7'h3d == _state_T_4[6:0] ? $signed(array_61) : $signed(_GEN_221); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_223 = 7'h3e == _state_T_4[6:0] ? $signed(array_62) : $signed(_GEN_222); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_224 = 7'h3f == _state_T_4[6:0] ? $signed(array_63) : $signed(_GEN_223); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_225 = 7'h40 == _state_T_4[6:0] ? $signed(array_64) : $signed(_GEN_224); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_226 = 7'h41 == _state_T_4[6:0] ? $signed(array_65) : $signed(_GEN_225); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_227 = 7'h42 == _state_T_4[6:0] ? $signed(array_66) : $signed(_GEN_226); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_228 = 7'h43 == _state_T_4[6:0] ? $signed(array_67) : $signed(_GEN_227); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_229 = 7'h44 == _state_T_4[6:0] ? $signed(array_68) : $signed(_GEN_228); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_230 = 7'h45 == _state_T_4[6:0] ? $signed(array_69) : $signed(_GEN_229); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_231 = 7'h46 == _state_T_4[6:0] ? $signed(array_70) : $signed(_GEN_230); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_232 = 7'h47 == _state_T_4[6:0] ? $signed(array_71) : $signed(_GEN_231); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_233 = 7'h48 == _state_T_4[6:0] ? $signed(array_72) : $signed(_GEN_232); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_234 = 7'h49 == _state_T_4[6:0] ? $signed(array_73) : $signed(_GEN_233); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_235 = 7'h4a == _state_T_4[6:0] ? $signed(array_74) : $signed(_GEN_234); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_236 = 7'h4b == _state_T_4[6:0] ? $signed(array_75) : $signed(_GEN_235); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_237 = 7'h4c == _state_T_4[6:0] ? $signed(array_76) : $signed(_GEN_236); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_238 = 7'h4d == _state_T_4[6:0] ? $signed(array_77) : $signed(_GEN_237); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_239 = 7'h4e == _state_T_4[6:0] ? $signed(array_78) : $signed(_GEN_238); // @[insertSort.scala 46:{64,64}]
  wire [31:0] _GEN_240 = 7'h4f == _state_T_4[6:0] ? $signed(array_79) : $signed(_GEN_239); // @[insertSort.scala 46:{64,64}]
  wire  _state_T_6 = $signed(_GEN_240) > $signed(key); // @[insertSort.scala 46:64]
  wire [2:0] _state_T_8 = $signed(j) > 32'sh0 & $signed(_GEN_240) > $signed(key) ? 3'h5 : 3'h7; // @[insertSort.scala 46:25]
  wire [31:0] _T_12 = $signed(j) + 32'sh1; // @[insertSort.scala 49:42]
  wire [31:0] _GEN_241 = 7'h0 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_1); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_242 = 7'h1 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_2); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_243 = 7'h2 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_3); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_244 = 7'h3 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_4); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_245 = 7'h4 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_5); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_246 = 7'h5 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_6); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_247 = 7'h6 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_7); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_248 = 7'h7 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_8); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_249 = 7'h8 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_9); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_250 = 7'h9 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_10); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_251 = 7'ha == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_11); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_252 = 7'hb == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_12); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_253 = 7'hc == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_13); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_254 = 7'hd == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_14); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_255 = 7'he == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_15); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_256 = 7'hf == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_16); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_257 = 7'h10 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_17); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_258 = 7'h11 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_18); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_259 = 7'h12 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_19); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_260 = 7'h13 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_20); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_261 = 7'h14 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_21); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_262 = 7'h15 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_22); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_263 = 7'h16 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_23); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_264 = 7'h17 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_24); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_265 = 7'h18 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_25); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_266 = 7'h19 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_26); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_267 = 7'h1a == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_27); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_268 = 7'h1b == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_28); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_269 = 7'h1c == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_29); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_270 = 7'h1d == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_30); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_271 = 7'h1e == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_31); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_272 = 7'h1f == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_32); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_273 = 7'h20 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_33); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_274 = 7'h21 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_34); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_275 = 7'h22 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_35); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_276 = 7'h23 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_36); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_277 = 7'h24 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_37); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_278 = 7'h25 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_38); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_279 = 7'h26 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_39); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_280 = 7'h27 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_40); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_281 = 7'h28 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_41); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_282 = 7'h29 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_42); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_283 = 7'h2a == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_43); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_284 = 7'h2b == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_44); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_285 = 7'h2c == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_45); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_286 = 7'h2d == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_46); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_287 = 7'h2e == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_47); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_288 = 7'h2f == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_48); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_289 = 7'h30 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_49); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_290 = 7'h31 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_50); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_291 = 7'h32 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_51); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_292 = 7'h33 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_52); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_293 = 7'h34 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_53); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_294 = 7'h35 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_54); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_295 = 7'h36 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_55); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_296 = 7'h37 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_56); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_297 = 7'h38 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_57); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_298 = 7'h39 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_58); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_299 = 7'h3a == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_59); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_300 = 7'h3b == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_60); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_301 = 7'h3c == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_61); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_302 = 7'h3d == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_62); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_303 = 7'h3e == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_63); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_304 = 7'h3f == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_64); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_305 = 7'h40 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_65); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_306 = 7'h41 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_66); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_307 = 7'h42 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_67); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_308 = 7'h43 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_68); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_309 = 7'h44 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_69); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_310 = 7'h45 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_70); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_311 = 7'h46 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_71); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_312 = 7'h47 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_72); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_313 = 7'h48 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_73); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_314 = 7'h49 == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_74); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_315 = 7'h4a == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_75); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_316 = 7'h4b == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_76); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_317 = 7'h4c == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_77); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_318 = 7'h4d == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_78); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_319 = 7'h4e == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_79); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _GEN_320 = 7'h4f == _T_12[6:0] ? $signed(_GEN_240) : $signed(_GEN_80); // @[insertSort.scala 49:{46,46}]
  wire [31:0] _j_T_5 = $signed(j) - 32'sh1; // @[insertSort.scala 53:20]
  wire [3:0] _state_T_14 = $signed(j) == 32'sh0 & _state_T_6 ? 4'h8 : 4'ha; // @[insertSort.scala 57:25]
  wire [31:0] _GEN_641 = 7'h0 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_1); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_642 = 7'h1 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_2); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_643 = 7'h2 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_3); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_644 = 7'h3 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_4); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_645 = 7'h4 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_5); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_646 = 7'h5 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_6); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_647 = 7'h6 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_7); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_648 = 7'h7 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_8); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_649 = 7'h8 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_9); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_650 = 7'h9 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_10); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_651 = 7'ha == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_11); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_652 = 7'hb == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_12); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_653 = 7'hc == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_13); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_654 = 7'hd == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_14); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_655 = 7'he == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_15); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_656 = 7'hf == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_16); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_657 = 7'h10 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_17); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_658 = 7'h11 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_18); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_659 = 7'h12 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_19); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_660 = 7'h13 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_20); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_661 = 7'h14 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_21); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_662 = 7'h15 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_22); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_663 = 7'h16 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_23); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_664 = 7'h17 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_24); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_665 = 7'h18 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_25); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_666 = 7'h19 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_26); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_667 = 7'h1a == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_27); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_668 = 7'h1b == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_28); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_669 = 7'h1c == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_29); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_670 = 7'h1d == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_30); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_671 = 7'h1e == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_31); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_672 = 7'h1f == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_32); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_673 = 7'h20 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_33); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_674 = 7'h21 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_34); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_675 = 7'h22 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_35); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_676 = 7'h23 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_36); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_677 = 7'h24 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_37); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_678 = 7'h25 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_38); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_679 = 7'h26 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_39); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_680 = 7'h27 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_40); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_681 = 7'h28 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_41); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_682 = 7'h29 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_42); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_683 = 7'h2a == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_43); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_684 = 7'h2b == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_44); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_685 = 7'h2c == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_45); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_686 = 7'h2d == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_46); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_687 = 7'h2e == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_47); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_688 = 7'h2f == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_48); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_689 = 7'h30 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_49); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_690 = 7'h31 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_50); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_691 = 7'h32 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_51); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_692 = 7'h33 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_52); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_693 = 7'h34 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_53); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_694 = 7'h35 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_54); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_695 = 7'h36 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_55); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_696 = 7'h37 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_56); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_697 = 7'h38 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_57); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_698 = 7'h39 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_58); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_699 = 7'h3a == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_59); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_700 = 7'h3b == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_60); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_701 = 7'h3c == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_61); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_702 = 7'h3d == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_62); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_703 = 7'h3e == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_63); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_704 = 7'h3f == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_64); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_705 = 7'h40 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_65); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_706 = 7'h41 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_66); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_707 = 7'h42 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_67); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_708 = 7'h43 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_68); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_709 = 7'h44 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_69); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_710 = 7'h45 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_70); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_711 = 7'h46 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_71); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_712 = 7'h47 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_72); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_713 = 7'h48 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_73); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_714 = 7'h49 == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_74); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_715 = 7'h4a == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_75); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_716 = 7'h4b == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_76); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_717 = 7'h4c == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_77); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_718 = 7'h4d == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_78); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_719 = 7'h4e == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_79); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_720 = 7'h4f == _state_T_4[6:0] ? $signed(key) : $signed(_GEN_80); // @[insertSort.scala 64:{33,33}]
  wire [31:0] _GEN_721 = 7'h0 == _T_12[6:0] ? $signed(key) : $signed(_GEN_1); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_722 = 7'h1 == _T_12[6:0] ? $signed(key) : $signed(_GEN_2); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_723 = 7'h2 == _T_12[6:0] ? $signed(key) : $signed(_GEN_3); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_724 = 7'h3 == _T_12[6:0] ? $signed(key) : $signed(_GEN_4); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_725 = 7'h4 == _T_12[6:0] ? $signed(key) : $signed(_GEN_5); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_726 = 7'h5 == _T_12[6:0] ? $signed(key) : $signed(_GEN_6); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_727 = 7'h6 == _T_12[6:0] ? $signed(key) : $signed(_GEN_7); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_728 = 7'h7 == _T_12[6:0] ? $signed(key) : $signed(_GEN_8); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_729 = 7'h8 == _T_12[6:0] ? $signed(key) : $signed(_GEN_9); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_730 = 7'h9 == _T_12[6:0] ? $signed(key) : $signed(_GEN_10); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_731 = 7'ha == _T_12[6:0] ? $signed(key) : $signed(_GEN_11); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_732 = 7'hb == _T_12[6:0] ? $signed(key) : $signed(_GEN_12); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_733 = 7'hc == _T_12[6:0] ? $signed(key) : $signed(_GEN_13); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_734 = 7'hd == _T_12[6:0] ? $signed(key) : $signed(_GEN_14); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_735 = 7'he == _T_12[6:0] ? $signed(key) : $signed(_GEN_15); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_736 = 7'hf == _T_12[6:0] ? $signed(key) : $signed(_GEN_16); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_737 = 7'h10 == _T_12[6:0] ? $signed(key) : $signed(_GEN_17); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_738 = 7'h11 == _T_12[6:0] ? $signed(key) : $signed(_GEN_18); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_739 = 7'h12 == _T_12[6:0] ? $signed(key) : $signed(_GEN_19); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_740 = 7'h13 == _T_12[6:0] ? $signed(key) : $signed(_GEN_20); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_741 = 7'h14 == _T_12[6:0] ? $signed(key) : $signed(_GEN_21); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_742 = 7'h15 == _T_12[6:0] ? $signed(key) : $signed(_GEN_22); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_743 = 7'h16 == _T_12[6:0] ? $signed(key) : $signed(_GEN_23); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_744 = 7'h17 == _T_12[6:0] ? $signed(key) : $signed(_GEN_24); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_745 = 7'h18 == _T_12[6:0] ? $signed(key) : $signed(_GEN_25); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_746 = 7'h19 == _T_12[6:0] ? $signed(key) : $signed(_GEN_26); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_747 = 7'h1a == _T_12[6:0] ? $signed(key) : $signed(_GEN_27); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_748 = 7'h1b == _T_12[6:0] ? $signed(key) : $signed(_GEN_28); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_749 = 7'h1c == _T_12[6:0] ? $signed(key) : $signed(_GEN_29); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_750 = 7'h1d == _T_12[6:0] ? $signed(key) : $signed(_GEN_30); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_751 = 7'h1e == _T_12[6:0] ? $signed(key) : $signed(_GEN_31); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_752 = 7'h1f == _T_12[6:0] ? $signed(key) : $signed(_GEN_32); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_753 = 7'h20 == _T_12[6:0] ? $signed(key) : $signed(_GEN_33); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_754 = 7'h21 == _T_12[6:0] ? $signed(key) : $signed(_GEN_34); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_755 = 7'h22 == _T_12[6:0] ? $signed(key) : $signed(_GEN_35); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_756 = 7'h23 == _T_12[6:0] ? $signed(key) : $signed(_GEN_36); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_757 = 7'h24 == _T_12[6:0] ? $signed(key) : $signed(_GEN_37); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_758 = 7'h25 == _T_12[6:0] ? $signed(key) : $signed(_GEN_38); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_759 = 7'h26 == _T_12[6:0] ? $signed(key) : $signed(_GEN_39); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_760 = 7'h27 == _T_12[6:0] ? $signed(key) : $signed(_GEN_40); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_761 = 7'h28 == _T_12[6:0] ? $signed(key) : $signed(_GEN_41); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_762 = 7'h29 == _T_12[6:0] ? $signed(key) : $signed(_GEN_42); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_763 = 7'h2a == _T_12[6:0] ? $signed(key) : $signed(_GEN_43); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_764 = 7'h2b == _T_12[6:0] ? $signed(key) : $signed(_GEN_44); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_765 = 7'h2c == _T_12[6:0] ? $signed(key) : $signed(_GEN_45); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_766 = 7'h2d == _T_12[6:0] ? $signed(key) : $signed(_GEN_46); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_767 = 7'h2e == _T_12[6:0] ? $signed(key) : $signed(_GEN_47); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_768 = 7'h2f == _T_12[6:0] ? $signed(key) : $signed(_GEN_48); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_769 = 7'h30 == _T_12[6:0] ? $signed(key) : $signed(_GEN_49); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_770 = 7'h31 == _T_12[6:0] ? $signed(key) : $signed(_GEN_50); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_771 = 7'h32 == _T_12[6:0] ? $signed(key) : $signed(_GEN_51); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_772 = 7'h33 == _T_12[6:0] ? $signed(key) : $signed(_GEN_52); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_773 = 7'h34 == _T_12[6:0] ? $signed(key) : $signed(_GEN_53); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_774 = 7'h35 == _T_12[6:0] ? $signed(key) : $signed(_GEN_54); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_775 = 7'h36 == _T_12[6:0] ? $signed(key) : $signed(_GEN_55); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_776 = 7'h37 == _T_12[6:0] ? $signed(key) : $signed(_GEN_56); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_777 = 7'h38 == _T_12[6:0] ? $signed(key) : $signed(_GEN_57); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_778 = 7'h39 == _T_12[6:0] ? $signed(key) : $signed(_GEN_58); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_779 = 7'h3a == _T_12[6:0] ? $signed(key) : $signed(_GEN_59); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_780 = 7'h3b == _T_12[6:0] ? $signed(key) : $signed(_GEN_60); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_781 = 7'h3c == _T_12[6:0] ? $signed(key) : $signed(_GEN_61); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_782 = 7'h3d == _T_12[6:0] ? $signed(key) : $signed(_GEN_62); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_783 = 7'h3e == _T_12[6:0] ? $signed(key) : $signed(_GEN_63); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_784 = 7'h3f == _T_12[6:0] ? $signed(key) : $signed(_GEN_64); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_785 = 7'h40 == _T_12[6:0] ? $signed(key) : $signed(_GEN_65); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_786 = 7'h41 == _T_12[6:0] ? $signed(key) : $signed(_GEN_66); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_787 = 7'h42 == _T_12[6:0] ? $signed(key) : $signed(_GEN_67); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_788 = 7'h43 == _T_12[6:0] ? $signed(key) : $signed(_GEN_68); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_789 = 7'h44 == _T_12[6:0] ? $signed(key) : $signed(_GEN_69); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_790 = 7'h45 == _T_12[6:0] ? $signed(key) : $signed(_GEN_70); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_791 = 7'h46 == _T_12[6:0] ? $signed(key) : $signed(_GEN_71); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_792 = 7'h47 == _T_12[6:0] ? $signed(key) : $signed(_GEN_72); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_793 = 7'h48 == _T_12[6:0] ? $signed(key) : $signed(_GEN_73); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_794 = 7'h49 == _T_12[6:0] ? $signed(key) : $signed(_GEN_74); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_795 = 7'h4a == _T_12[6:0] ? $signed(key) : $signed(_GEN_75); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_796 = 7'h4b == _T_12[6:0] ? $signed(key) : $signed(_GEN_76); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_797 = 7'h4c == _T_12[6:0] ? $signed(key) : $signed(_GEN_77); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_798 = 7'h4d == _T_12[6:0] ? $signed(key) : $signed(_GEN_78); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_799 = 7'h4e == _T_12[6:0] ? $signed(key) : $signed(_GEN_79); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _GEN_800 = 7'h4f == _T_12[6:0] ? $signed(key) : $signed(_GEN_80); // @[insertSort.scala 68:{46,46}]
  wire [31:0] _i_T_2 = $signed(i) + 32'sh1; // @[insertSort.scala 72:21]
  wire [3:0] _GEN_801 = 4'hc == state ? 4'hf : _GEN_0; // @[insertSort.scala 26:19 76:19]
  wire [31:0] _GEN_802 = 4'hb == state ? $signed(_i_T_2) : $signed(i); // @[insertSort.scala 26:19 72:15 22:16]
  wire [3:0] _GEN_803 = 4'hb == state ? 4'h1 : _GEN_801; // @[insertSort.scala 26:19 73:19]
  wire [31:0] _GEN_804 = 4'ha == state ? $signed(_GEN_721) : $signed(_GEN_1); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_805 = 4'ha == state ? $signed(_GEN_722) : $signed(_GEN_2); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_806 = 4'ha == state ? $signed(_GEN_723) : $signed(_GEN_3); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_807 = 4'ha == state ? $signed(_GEN_724) : $signed(_GEN_4); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_808 = 4'ha == state ? $signed(_GEN_725) : $signed(_GEN_5); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_809 = 4'ha == state ? $signed(_GEN_726) : $signed(_GEN_6); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_810 = 4'ha == state ? $signed(_GEN_727) : $signed(_GEN_7); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_811 = 4'ha == state ? $signed(_GEN_728) : $signed(_GEN_8); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_812 = 4'ha == state ? $signed(_GEN_729) : $signed(_GEN_9); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_813 = 4'ha == state ? $signed(_GEN_730) : $signed(_GEN_10); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_814 = 4'ha == state ? $signed(_GEN_731) : $signed(_GEN_11); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_815 = 4'ha == state ? $signed(_GEN_732) : $signed(_GEN_12); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_816 = 4'ha == state ? $signed(_GEN_733) : $signed(_GEN_13); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_817 = 4'ha == state ? $signed(_GEN_734) : $signed(_GEN_14); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_818 = 4'ha == state ? $signed(_GEN_735) : $signed(_GEN_15); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_819 = 4'ha == state ? $signed(_GEN_736) : $signed(_GEN_16); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_820 = 4'ha == state ? $signed(_GEN_737) : $signed(_GEN_17); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_821 = 4'ha == state ? $signed(_GEN_738) : $signed(_GEN_18); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_822 = 4'ha == state ? $signed(_GEN_739) : $signed(_GEN_19); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_823 = 4'ha == state ? $signed(_GEN_740) : $signed(_GEN_20); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_824 = 4'ha == state ? $signed(_GEN_741) : $signed(_GEN_21); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_825 = 4'ha == state ? $signed(_GEN_742) : $signed(_GEN_22); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_826 = 4'ha == state ? $signed(_GEN_743) : $signed(_GEN_23); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_827 = 4'ha == state ? $signed(_GEN_744) : $signed(_GEN_24); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_828 = 4'ha == state ? $signed(_GEN_745) : $signed(_GEN_25); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_829 = 4'ha == state ? $signed(_GEN_746) : $signed(_GEN_26); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_830 = 4'ha == state ? $signed(_GEN_747) : $signed(_GEN_27); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_831 = 4'ha == state ? $signed(_GEN_748) : $signed(_GEN_28); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_832 = 4'ha == state ? $signed(_GEN_749) : $signed(_GEN_29); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_833 = 4'ha == state ? $signed(_GEN_750) : $signed(_GEN_30); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_834 = 4'ha == state ? $signed(_GEN_751) : $signed(_GEN_31); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_835 = 4'ha == state ? $signed(_GEN_752) : $signed(_GEN_32); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_836 = 4'ha == state ? $signed(_GEN_753) : $signed(_GEN_33); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_837 = 4'ha == state ? $signed(_GEN_754) : $signed(_GEN_34); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_838 = 4'ha == state ? $signed(_GEN_755) : $signed(_GEN_35); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_839 = 4'ha == state ? $signed(_GEN_756) : $signed(_GEN_36); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_840 = 4'ha == state ? $signed(_GEN_757) : $signed(_GEN_37); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_841 = 4'ha == state ? $signed(_GEN_758) : $signed(_GEN_38); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_842 = 4'ha == state ? $signed(_GEN_759) : $signed(_GEN_39); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_843 = 4'ha == state ? $signed(_GEN_760) : $signed(_GEN_40); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_844 = 4'ha == state ? $signed(_GEN_761) : $signed(_GEN_41); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_845 = 4'ha == state ? $signed(_GEN_762) : $signed(_GEN_42); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_846 = 4'ha == state ? $signed(_GEN_763) : $signed(_GEN_43); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_847 = 4'ha == state ? $signed(_GEN_764) : $signed(_GEN_44); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_848 = 4'ha == state ? $signed(_GEN_765) : $signed(_GEN_45); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_849 = 4'ha == state ? $signed(_GEN_766) : $signed(_GEN_46); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_850 = 4'ha == state ? $signed(_GEN_767) : $signed(_GEN_47); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_851 = 4'ha == state ? $signed(_GEN_768) : $signed(_GEN_48); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_852 = 4'ha == state ? $signed(_GEN_769) : $signed(_GEN_49); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_853 = 4'ha == state ? $signed(_GEN_770) : $signed(_GEN_50); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_854 = 4'ha == state ? $signed(_GEN_771) : $signed(_GEN_51); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_855 = 4'ha == state ? $signed(_GEN_772) : $signed(_GEN_52); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_856 = 4'ha == state ? $signed(_GEN_773) : $signed(_GEN_53); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_857 = 4'ha == state ? $signed(_GEN_774) : $signed(_GEN_54); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_858 = 4'ha == state ? $signed(_GEN_775) : $signed(_GEN_55); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_859 = 4'ha == state ? $signed(_GEN_776) : $signed(_GEN_56); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_860 = 4'ha == state ? $signed(_GEN_777) : $signed(_GEN_57); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_861 = 4'ha == state ? $signed(_GEN_778) : $signed(_GEN_58); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_862 = 4'ha == state ? $signed(_GEN_779) : $signed(_GEN_59); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_863 = 4'ha == state ? $signed(_GEN_780) : $signed(_GEN_60); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_864 = 4'ha == state ? $signed(_GEN_781) : $signed(_GEN_61); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_865 = 4'ha == state ? $signed(_GEN_782) : $signed(_GEN_62); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_866 = 4'ha == state ? $signed(_GEN_783) : $signed(_GEN_63); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_867 = 4'ha == state ? $signed(_GEN_784) : $signed(_GEN_64); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_868 = 4'ha == state ? $signed(_GEN_785) : $signed(_GEN_65); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_869 = 4'ha == state ? $signed(_GEN_786) : $signed(_GEN_66); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_870 = 4'ha == state ? $signed(_GEN_787) : $signed(_GEN_67); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_871 = 4'ha == state ? $signed(_GEN_788) : $signed(_GEN_68); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_872 = 4'ha == state ? $signed(_GEN_789) : $signed(_GEN_69); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_873 = 4'ha == state ? $signed(_GEN_790) : $signed(_GEN_70); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_874 = 4'ha == state ? $signed(_GEN_791) : $signed(_GEN_71); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_875 = 4'ha == state ? $signed(_GEN_792) : $signed(_GEN_72); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_876 = 4'ha == state ? $signed(_GEN_793) : $signed(_GEN_73); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_877 = 4'ha == state ? $signed(_GEN_794) : $signed(_GEN_74); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_878 = 4'ha == state ? $signed(_GEN_795) : $signed(_GEN_75); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_879 = 4'ha == state ? $signed(_GEN_796) : $signed(_GEN_76); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_880 = 4'ha == state ? $signed(_GEN_797) : $signed(_GEN_77); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_881 = 4'ha == state ? $signed(_GEN_798) : $signed(_GEN_78); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_882 = 4'ha == state ? $signed(_GEN_799) : $signed(_GEN_79); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_883 = 4'ha == state ? $signed(_GEN_800) : $signed(_GEN_80); // @[insertSort.scala 26:19]
  wire [3:0] _GEN_884 = 4'ha == state ? 4'hb : _GEN_803; // @[insertSort.scala 26:19 69:19]
  wire [31:0] _GEN_885 = 4'ha == state ? $signed(i) : $signed(_GEN_802); // @[insertSort.scala 22:16 26:19]
  wire [31:0] _GEN_886 = 4'h9 == state ? $signed(_GEN_641) : $signed(_GEN_804); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_887 = 4'h9 == state ? $signed(_GEN_642) : $signed(_GEN_805); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_888 = 4'h9 == state ? $signed(_GEN_643) : $signed(_GEN_806); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_889 = 4'h9 == state ? $signed(_GEN_644) : $signed(_GEN_807); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_890 = 4'h9 == state ? $signed(_GEN_645) : $signed(_GEN_808); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_891 = 4'h9 == state ? $signed(_GEN_646) : $signed(_GEN_809); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_892 = 4'h9 == state ? $signed(_GEN_647) : $signed(_GEN_810); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_893 = 4'h9 == state ? $signed(_GEN_648) : $signed(_GEN_811); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_894 = 4'h9 == state ? $signed(_GEN_649) : $signed(_GEN_812); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_895 = 4'h9 == state ? $signed(_GEN_650) : $signed(_GEN_813); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_896 = 4'h9 == state ? $signed(_GEN_651) : $signed(_GEN_814); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_897 = 4'h9 == state ? $signed(_GEN_652) : $signed(_GEN_815); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_898 = 4'h9 == state ? $signed(_GEN_653) : $signed(_GEN_816); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_899 = 4'h9 == state ? $signed(_GEN_654) : $signed(_GEN_817); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_900 = 4'h9 == state ? $signed(_GEN_655) : $signed(_GEN_818); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_901 = 4'h9 == state ? $signed(_GEN_656) : $signed(_GEN_819); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_902 = 4'h9 == state ? $signed(_GEN_657) : $signed(_GEN_820); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_903 = 4'h9 == state ? $signed(_GEN_658) : $signed(_GEN_821); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_904 = 4'h9 == state ? $signed(_GEN_659) : $signed(_GEN_822); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_905 = 4'h9 == state ? $signed(_GEN_660) : $signed(_GEN_823); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_906 = 4'h9 == state ? $signed(_GEN_661) : $signed(_GEN_824); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_907 = 4'h9 == state ? $signed(_GEN_662) : $signed(_GEN_825); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_908 = 4'h9 == state ? $signed(_GEN_663) : $signed(_GEN_826); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_909 = 4'h9 == state ? $signed(_GEN_664) : $signed(_GEN_827); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_910 = 4'h9 == state ? $signed(_GEN_665) : $signed(_GEN_828); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_911 = 4'h9 == state ? $signed(_GEN_666) : $signed(_GEN_829); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_912 = 4'h9 == state ? $signed(_GEN_667) : $signed(_GEN_830); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_913 = 4'h9 == state ? $signed(_GEN_668) : $signed(_GEN_831); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_914 = 4'h9 == state ? $signed(_GEN_669) : $signed(_GEN_832); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_915 = 4'h9 == state ? $signed(_GEN_670) : $signed(_GEN_833); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_916 = 4'h9 == state ? $signed(_GEN_671) : $signed(_GEN_834); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_917 = 4'h9 == state ? $signed(_GEN_672) : $signed(_GEN_835); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_918 = 4'h9 == state ? $signed(_GEN_673) : $signed(_GEN_836); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_919 = 4'h9 == state ? $signed(_GEN_674) : $signed(_GEN_837); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_920 = 4'h9 == state ? $signed(_GEN_675) : $signed(_GEN_838); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_921 = 4'h9 == state ? $signed(_GEN_676) : $signed(_GEN_839); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_922 = 4'h9 == state ? $signed(_GEN_677) : $signed(_GEN_840); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_923 = 4'h9 == state ? $signed(_GEN_678) : $signed(_GEN_841); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_924 = 4'h9 == state ? $signed(_GEN_679) : $signed(_GEN_842); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_925 = 4'h9 == state ? $signed(_GEN_680) : $signed(_GEN_843); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_926 = 4'h9 == state ? $signed(_GEN_681) : $signed(_GEN_844); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_927 = 4'h9 == state ? $signed(_GEN_682) : $signed(_GEN_845); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_928 = 4'h9 == state ? $signed(_GEN_683) : $signed(_GEN_846); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_929 = 4'h9 == state ? $signed(_GEN_684) : $signed(_GEN_847); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_930 = 4'h9 == state ? $signed(_GEN_685) : $signed(_GEN_848); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_931 = 4'h9 == state ? $signed(_GEN_686) : $signed(_GEN_849); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_932 = 4'h9 == state ? $signed(_GEN_687) : $signed(_GEN_850); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_933 = 4'h9 == state ? $signed(_GEN_688) : $signed(_GEN_851); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_934 = 4'h9 == state ? $signed(_GEN_689) : $signed(_GEN_852); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_935 = 4'h9 == state ? $signed(_GEN_690) : $signed(_GEN_853); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_936 = 4'h9 == state ? $signed(_GEN_691) : $signed(_GEN_854); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_937 = 4'h9 == state ? $signed(_GEN_692) : $signed(_GEN_855); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_938 = 4'h9 == state ? $signed(_GEN_693) : $signed(_GEN_856); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_939 = 4'h9 == state ? $signed(_GEN_694) : $signed(_GEN_857); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_940 = 4'h9 == state ? $signed(_GEN_695) : $signed(_GEN_858); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_941 = 4'h9 == state ? $signed(_GEN_696) : $signed(_GEN_859); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_942 = 4'h9 == state ? $signed(_GEN_697) : $signed(_GEN_860); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_943 = 4'h9 == state ? $signed(_GEN_698) : $signed(_GEN_861); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_944 = 4'h9 == state ? $signed(_GEN_699) : $signed(_GEN_862); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_945 = 4'h9 == state ? $signed(_GEN_700) : $signed(_GEN_863); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_946 = 4'h9 == state ? $signed(_GEN_701) : $signed(_GEN_864); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_947 = 4'h9 == state ? $signed(_GEN_702) : $signed(_GEN_865); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_948 = 4'h9 == state ? $signed(_GEN_703) : $signed(_GEN_866); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_949 = 4'h9 == state ? $signed(_GEN_704) : $signed(_GEN_867); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_950 = 4'h9 == state ? $signed(_GEN_705) : $signed(_GEN_868); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_951 = 4'h9 == state ? $signed(_GEN_706) : $signed(_GEN_869); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_952 = 4'h9 == state ? $signed(_GEN_707) : $signed(_GEN_870); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_953 = 4'h9 == state ? $signed(_GEN_708) : $signed(_GEN_871); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_954 = 4'h9 == state ? $signed(_GEN_709) : $signed(_GEN_872); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_955 = 4'h9 == state ? $signed(_GEN_710) : $signed(_GEN_873); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_956 = 4'h9 == state ? $signed(_GEN_711) : $signed(_GEN_874); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_957 = 4'h9 == state ? $signed(_GEN_712) : $signed(_GEN_875); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_958 = 4'h9 == state ? $signed(_GEN_713) : $signed(_GEN_876); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_959 = 4'h9 == state ? $signed(_GEN_714) : $signed(_GEN_877); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_960 = 4'h9 == state ? $signed(_GEN_715) : $signed(_GEN_878); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_961 = 4'h9 == state ? $signed(_GEN_716) : $signed(_GEN_879); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_962 = 4'h9 == state ? $signed(_GEN_717) : $signed(_GEN_880); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_963 = 4'h9 == state ? $signed(_GEN_718) : $signed(_GEN_881); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_964 = 4'h9 == state ? $signed(_GEN_719) : $signed(_GEN_882); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_965 = 4'h9 == state ? $signed(_GEN_720) : $signed(_GEN_883); // @[insertSort.scala 26:19]
  wire [3:0] _GEN_966 = 4'h9 == state ? 4'hb : _GEN_884; // @[insertSort.scala 26:19 65:19]
  wire [31:0] _GEN_967 = 4'h9 == state ? $signed(i) : $signed(_GEN_885); // @[insertSort.scala 22:16 26:19]
  wire [31:0] _GEN_968 = 4'h8 == state ? $signed(_GEN_241) : $signed(_GEN_886); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_969 = 4'h8 == state ? $signed(_GEN_242) : $signed(_GEN_887); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_970 = 4'h8 == state ? $signed(_GEN_243) : $signed(_GEN_888); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_971 = 4'h8 == state ? $signed(_GEN_244) : $signed(_GEN_889); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_972 = 4'h8 == state ? $signed(_GEN_245) : $signed(_GEN_890); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_973 = 4'h8 == state ? $signed(_GEN_246) : $signed(_GEN_891); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_974 = 4'h8 == state ? $signed(_GEN_247) : $signed(_GEN_892); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_975 = 4'h8 == state ? $signed(_GEN_248) : $signed(_GEN_893); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_976 = 4'h8 == state ? $signed(_GEN_249) : $signed(_GEN_894); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_977 = 4'h8 == state ? $signed(_GEN_250) : $signed(_GEN_895); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_978 = 4'h8 == state ? $signed(_GEN_251) : $signed(_GEN_896); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_979 = 4'h8 == state ? $signed(_GEN_252) : $signed(_GEN_897); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_980 = 4'h8 == state ? $signed(_GEN_253) : $signed(_GEN_898); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_981 = 4'h8 == state ? $signed(_GEN_254) : $signed(_GEN_899); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_982 = 4'h8 == state ? $signed(_GEN_255) : $signed(_GEN_900); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_983 = 4'h8 == state ? $signed(_GEN_256) : $signed(_GEN_901); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_984 = 4'h8 == state ? $signed(_GEN_257) : $signed(_GEN_902); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_985 = 4'h8 == state ? $signed(_GEN_258) : $signed(_GEN_903); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_986 = 4'h8 == state ? $signed(_GEN_259) : $signed(_GEN_904); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_987 = 4'h8 == state ? $signed(_GEN_260) : $signed(_GEN_905); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_988 = 4'h8 == state ? $signed(_GEN_261) : $signed(_GEN_906); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_989 = 4'h8 == state ? $signed(_GEN_262) : $signed(_GEN_907); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_990 = 4'h8 == state ? $signed(_GEN_263) : $signed(_GEN_908); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_991 = 4'h8 == state ? $signed(_GEN_264) : $signed(_GEN_909); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_992 = 4'h8 == state ? $signed(_GEN_265) : $signed(_GEN_910); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_993 = 4'h8 == state ? $signed(_GEN_266) : $signed(_GEN_911); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_994 = 4'h8 == state ? $signed(_GEN_267) : $signed(_GEN_912); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_995 = 4'h8 == state ? $signed(_GEN_268) : $signed(_GEN_913); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_996 = 4'h8 == state ? $signed(_GEN_269) : $signed(_GEN_914); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_997 = 4'h8 == state ? $signed(_GEN_270) : $signed(_GEN_915); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_998 = 4'h8 == state ? $signed(_GEN_271) : $signed(_GEN_916); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_999 = 4'h8 == state ? $signed(_GEN_272) : $signed(_GEN_917); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1000 = 4'h8 == state ? $signed(_GEN_273) : $signed(_GEN_918); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1001 = 4'h8 == state ? $signed(_GEN_274) : $signed(_GEN_919); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1002 = 4'h8 == state ? $signed(_GEN_275) : $signed(_GEN_920); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1003 = 4'h8 == state ? $signed(_GEN_276) : $signed(_GEN_921); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1004 = 4'h8 == state ? $signed(_GEN_277) : $signed(_GEN_922); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1005 = 4'h8 == state ? $signed(_GEN_278) : $signed(_GEN_923); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1006 = 4'h8 == state ? $signed(_GEN_279) : $signed(_GEN_924); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1007 = 4'h8 == state ? $signed(_GEN_280) : $signed(_GEN_925); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1008 = 4'h8 == state ? $signed(_GEN_281) : $signed(_GEN_926); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1009 = 4'h8 == state ? $signed(_GEN_282) : $signed(_GEN_927); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1010 = 4'h8 == state ? $signed(_GEN_283) : $signed(_GEN_928); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1011 = 4'h8 == state ? $signed(_GEN_284) : $signed(_GEN_929); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1012 = 4'h8 == state ? $signed(_GEN_285) : $signed(_GEN_930); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1013 = 4'h8 == state ? $signed(_GEN_286) : $signed(_GEN_931); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1014 = 4'h8 == state ? $signed(_GEN_287) : $signed(_GEN_932); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1015 = 4'h8 == state ? $signed(_GEN_288) : $signed(_GEN_933); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1016 = 4'h8 == state ? $signed(_GEN_289) : $signed(_GEN_934); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1017 = 4'h8 == state ? $signed(_GEN_290) : $signed(_GEN_935); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1018 = 4'h8 == state ? $signed(_GEN_291) : $signed(_GEN_936); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1019 = 4'h8 == state ? $signed(_GEN_292) : $signed(_GEN_937); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1020 = 4'h8 == state ? $signed(_GEN_293) : $signed(_GEN_938); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1021 = 4'h8 == state ? $signed(_GEN_294) : $signed(_GEN_939); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1022 = 4'h8 == state ? $signed(_GEN_295) : $signed(_GEN_940); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1023 = 4'h8 == state ? $signed(_GEN_296) : $signed(_GEN_941); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1024 = 4'h8 == state ? $signed(_GEN_297) : $signed(_GEN_942); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1025 = 4'h8 == state ? $signed(_GEN_298) : $signed(_GEN_943); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1026 = 4'h8 == state ? $signed(_GEN_299) : $signed(_GEN_944); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1027 = 4'h8 == state ? $signed(_GEN_300) : $signed(_GEN_945); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1028 = 4'h8 == state ? $signed(_GEN_301) : $signed(_GEN_946); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1029 = 4'h8 == state ? $signed(_GEN_302) : $signed(_GEN_947); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1030 = 4'h8 == state ? $signed(_GEN_303) : $signed(_GEN_948); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1031 = 4'h8 == state ? $signed(_GEN_304) : $signed(_GEN_949); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1032 = 4'h8 == state ? $signed(_GEN_305) : $signed(_GEN_950); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1033 = 4'h8 == state ? $signed(_GEN_306) : $signed(_GEN_951); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1034 = 4'h8 == state ? $signed(_GEN_307) : $signed(_GEN_952); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1035 = 4'h8 == state ? $signed(_GEN_308) : $signed(_GEN_953); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1036 = 4'h8 == state ? $signed(_GEN_309) : $signed(_GEN_954); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1037 = 4'h8 == state ? $signed(_GEN_310) : $signed(_GEN_955); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1038 = 4'h8 == state ? $signed(_GEN_311) : $signed(_GEN_956); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1039 = 4'h8 == state ? $signed(_GEN_312) : $signed(_GEN_957); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1040 = 4'h8 == state ? $signed(_GEN_313) : $signed(_GEN_958); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1041 = 4'h8 == state ? $signed(_GEN_314) : $signed(_GEN_959); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1042 = 4'h8 == state ? $signed(_GEN_315) : $signed(_GEN_960); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1043 = 4'h8 == state ? $signed(_GEN_316) : $signed(_GEN_961); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1044 = 4'h8 == state ? $signed(_GEN_317) : $signed(_GEN_962); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1045 = 4'h8 == state ? $signed(_GEN_318) : $signed(_GEN_963); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1046 = 4'h8 == state ? $signed(_GEN_319) : $signed(_GEN_964); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1047 = 4'h8 == state ? $signed(_GEN_320) : $signed(_GEN_965); // @[insertSort.scala 26:19]
  wire [3:0] _GEN_1048 = 4'h8 == state ? 4'h9 : _GEN_966; // @[insertSort.scala 26:19 61:19]
  wire [31:0] _GEN_1049 = 4'h8 == state ? $signed(i) : $signed(_GEN_967); // @[insertSort.scala 22:16 26:19]
  wire [3:0] _GEN_1050 = 4'h7 == state ? _state_T_14 : _GEN_1048; // @[insertSort.scala 26:19 57:19]
  wire [31:0] _GEN_1051 = 4'h7 == state ? $signed(_GEN_1) : $signed(_GEN_968); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1052 = 4'h7 == state ? $signed(_GEN_2) : $signed(_GEN_969); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1053 = 4'h7 == state ? $signed(_GEN_3) : $signed(_GEN_970); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1054 = 4'h7 == state ? $signed(_GEN_4) : $signed(_GEN_971); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1055 = 4'h7 == state ? $signed(_GEN_5) : $signed(_GEN_972); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1056 = 4'h7 == state ? $signed(_GEN_6) : $signed(_GEN_973); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1057 = 4'h7 == state ? $signed(_GEN_7) : $signed(_GEN_974); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1058 = 4'h7 == state ? $signed(_GEN_8) : $signed(_GEN_975); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1059 = 4'h7 == state ? $signed(_GEN_9) : $signed(_GEN_976); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1060 = 4'h7 == state ? $signed(_GEN_10) : $signed(_GEN_977); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1061 = 4'h7 == state ? $signed(_GEN_11) : $signed(_GEN_978); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1062 = 4'h7 == state ? $signed(_GEN_12) : $signed(_GEN_979); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1063 = 4'h7 == state ? $signed(_GEN_13) : $signed(_GEN_980); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1064 = 4'h7 == state ? $signed(_GEN_14) : $signed(_GEN_981); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1065 = 4'h7 == state ? $signed(_GEN_15) : $signed(_GEN_982); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1066 = 4'h7 == state ? $signed(_GEN_16) : $signed(_GEN_983); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1067 = 4'h7 == state ? $signed(_GEN_17) : $signed(_GEN_984); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1068 = 4'h7 == state ? $signed(_GEN_18) : $signed(_GEN_985); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1069 = 4'h7 == state ? $signed(_GEN_19) : $signed(_GEN_986); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1070 = 4'h7 == state ? $signed(_GEN_20) : $signed(_GEN_987); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1071 = 4'h7 == state ? $signed(_GEN_21) : $signed(_GEN_988); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1072 = 4'h7 == state ? $signed(_GEN_22) : $signed(_GEN_989); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1073 = 4'h7 == state ? $signed(_GEN_23) : $signed(_GEN_990); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1074 = 4'h7 == state ? $signed(_GEN_24) : $signed(_GEN_991); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1075 = 4'h7 == state ? $signed(_GEN_25) : $signed(_GEN_992); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1076 = 4'h7 == state ? $signed(_GEN_26) : $signed(_GEN_993); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1077 = 4'h7 == state ? $signed(_GEN_27) : $signed(_GEN_994); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1078 = 4'h7 == state ? $signed(_GEN_28) : $signed(_GEN_995); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1079 = 4'h7 == state ? $signed(_GEN_29) : $signed(_GEN_996); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1080 = 4'h7 == state ? $signed(_GEN_30) : $signed(_GEN_997); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1081 = 4'h7 == state ? $signed(_GEN_31) : $signed(_GEN_998); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1082 = 4'h7 == state ? $signed(_GEN_32) : $signed(_GEN_999); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1083 = 4'h7 == state ? $signed(_GEN_33) : $signed(_GEN_1000); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1084 = 4'h7 == state ? $signed(_GEN_34) : $signed(_GEN_1001); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1085 = 4'h7 == state ? $signed(_GEN_35) : $signed(_GEN_1002); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1086 = 4'h7 == state ? $signed(_GEN_36) : $signed(_GEN_1003); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1087 = 4'h7 == state ? $signed(_GEN_37) : $signed(_GEN_1004); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1088 = 4'h7 == state ? $signed(_GEN_38) : $signed(_GEN_1005); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1089 = 4'h7 == state ? $signed(_GEN_39) : $signed(_GEN_1006); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1090 = 4'h7 == state ? $signed(_GEN_40) : $signed(_GEN_1007); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1091 = 4'h7 == state ? $signed(_GEN_41) : $signed(_GEN_1008); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1092 = 4'h7 == state ? $signed(_GEN_42) : $signed(_GEN_1009); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1093 = 4'h7 == state ? $signed(_GEN_43) : $signed(_GEN_1010); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1094 = 4'h7 == state ? $signed(_GEN_44) : $signed(_GEN_1011); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1095 = 4'h7 == state ? $signed(_GEN_45) : $signed(_GEN_1012); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1096 = 4'h7 == state ? $signed(_GEN_46) : $signed(_GEN_1013); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1097 = 4'h7 == state ? $signed(_GEN_47) : $signed(_GEN_1014); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1098 = 4'h7 == state ? $signed(_GEN_48) : $signed(_GEN_1015); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1099 = 4'h7 == state ? $signed(_GEN_49) : $signed(_GEN_1016); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1100 = 4'h7 == state ? $signed(_GEN_50) : $signed(_GEN_1017); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1101 = 4'h7 == state ? $signed(_GEN_51) : $signed(_GEN_1018); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1102 = 4'h7 == state ? $signed(_GEN_52) : $signed(_GEN_1019); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1103 = 4'h7 == state ? $signed(_GEN_53) : $signed(_GEN_1020); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1104 = 4'h7 == state ? $signed(_GEN_54) : $signed(_GEN_1021); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1105 = 4'h7 == state ? $signed(_GEN_55) : $signed(_GEN_1022); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1106 = 4'h7 == state ? $signed(_GEN_56) : $signed(_GEN_1023); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1107 = 4'h7 == state ? $signed(_GEN_57) : $signed(_GEN_1024); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1108 = 4'h7 == state ? $signed(_GEN_58) : $signed(_GEN_1025); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1109 = 4'h7 == state ? $signed(_GEN_59) : $signed(_GEN_1026); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1110 = 4'h7 == state ? $signed(_GEN_60) : $signed(_GEN_1027); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1111 = 4'h7 == state ? $signed(_GEN_61) : $signed(_GEN_1028); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1112 = 4'h7 == state ? $signed(_GEN_62) : $signed(_GEN_1029); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1113 = 4'h7 == state ? $signed(_GEN_63) : $signed(_GEN_1030); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1114 = 4'h7 == state ? $signed(_GEN_64) : $signed(_GEN_1031); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1115 = 4'h7 == state ? $signed(_GEN_65) : $signed(_GEN_1032); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1116 = 4'h7 == state ? $signed(_GEN_66) : $signed(_GEN_1033); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1117 = 4'h7 == state ? $signed(_GEN_67) : $signed(_GEN_1034); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1118 = 4'h7 == state ? $signed(_GEN_68) : $signed(_GEN_1035); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1119 = 4'h7 == state ? $signed(_GEN_69) : $signed(_GEN_1036); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1120 = 4'h7 == state ? $signed(_GEN_70) : $signed(_GEN_1037); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1121 = 4'h7 == state ? $signed(_GEN_71) : $signed(_GEN_1038); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1122 = 4'h7 == state ? $signed(_GEN_72) : $signed(_GEN_1039); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1123 = 4'h7 == state ? $signed(_GEN_73) : $signed(_GEN_1040); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1124 = 4'h7 == state ? $signed(_GEN_74) : $signed(_GEN_1041); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1125 = 4'h7 == state ? $signed(_GEN_75) : $signed(_GEN_1042); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1126 = 4'h7 == state ? $signed(_GEN_76) : $signed(_GEN_1043); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1127 = 4'h7 == state ? $signed(_GEN_77) : $signed(_GEN_1044); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1128 = 4'h7 == state ? $signed(_GEN_78) : $signed(_GEN_1045); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1129 = 4'h7 == state ? $signed(_GEN_79) : $signed(_GEN_1046); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1130 = 4'h7 == state ? $signed(_GEN_80) : $signed(_GEN_1047); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1131 = 4'h7 == state ? $signed(i) : $signed(_GEN_1049); // @[insertSort.scala 22:16 26:19]
  wire [31:0] _GEN_1132 = 4'h6 == state ? $signed(_j_T_5) : $signed(j); // @[insertSort.scala 26:19 53:15 24:16]
  wire [3:0] _GEN_1133 = 4'h6 == state ? 4'h4 : _GEN_1050; // @[insertSort.scala 26:19 54:19]
  wire [31:0] _GEN_1134 = 4'h6 == state ? $signed(_GEN_1) : $signed(_GEN_1051); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1135 = 4'h6 == state ? $signed(_GEN_2) : $signed(_GEN_1052); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1136 = 4'h6 == state ? $signed(_GEN_3) : $signed(_GEN_1053); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1137 = 4'h6 == state ? $signed(_GEN_4) : $signed(_GEN_1054); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1138 = 4'h6 == state ? $signed(_GEN_5) : $signed(_GEN_1055); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1139 = 4'h6 == state ? $signed(_GEN_6) : $signed(_GEN_1056); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1140 = 4'h6 == state ? $signed(_GEN_7) : $signed(_GEN_1057); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1141 = 4'h6 == state ? $signed(_GEN_8) : $signed(_GEN_1058); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1142 = 4'h6 == state ? $signed(_GEN_9) : $signed(_GEN_1059); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1143 = 4'h6 == state ? $signed(_GEN_10) : $signed(_GEN_1060); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1144 = 4'h6 == state ? $signed(_GEN_11) : $signed(_GEN_1061); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1145 = 4'h6 == state ? $signed(_GEN_12) : $signed(_GEN_1062); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1146 = 4'h6 == state ? $signed(_GEN_13) : $signed(_GEN_1063); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1147 = 4'h6 == state ? $signed(_GEN_14) : $signed(_GEN_1064); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1148 = 4'h6 == state ? $signed(_GEN_15) : $signed(_GEN_1065); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1149 = 4'h6 == state ? $signed(_GEN_16) : $signed(_GEN_1066); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1150 = 4'h6 == state ? $signed(_GEN_17) : $signed(_GEN_1067); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1151 = 4'h6 == state ? $signed(_GEN_18) : $signed(_GEN_1068); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1152 = 4'h6 == state ? $signed(_GEN_19) : $signed(_GEN_1069); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1153 = 4'h6 == state ? $signed(_GEN_20) : $signed(_GEN_1070); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1154 = 4'h6 == state ? $signed(_GEN_21) : $signed(_GEN_1071); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1155 = 4'h6 == state ? $signed(_GEN_22) : $signed(_GEN_1072); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1156 = 4'h6 == state ? $signed(_GEN_23) : $signed(_GEN_1073); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1157 = 4'h6 == state ? $signed(_GEN_24) : $signed(_GEN_1074); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1158 = 4'h6 == state ? $signed(_GEN_25) : $signed(_GEN_1075); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1159 = 4'h6 == state ? $signed(_GEN_26) : $signed(_GEN_1076); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1160 = 4'h6 == state ? $signed(_GEN_27) : $signed(_GEN_1077); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1161 = 4'h6 == state ? $signed(_GEN_28) : $signed(_GEN_1078); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1162 = 4'h6 == state ? $signed(_GEN_29) : $signed(_GEN_1079); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1163 = 4'h6 == state ? $signed(_GEN_30) : $signed(_GEN_1080); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1164 = 4'h6 == state ? $signed(_GEN_31) : $signed(_GEN_1081); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1165 = 4'h6 == state ? $signed(_GEN_32) : $signed(_GEN_1082); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1166 = 4'h6 == state ? $signed(_GEN_33) : $signed(_GEN_1083); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1167 = 4'h6 == state ? $signed(_GEN_34) : $signed(_GEN_1084); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1168 = 4'h6 == state ? $signed(_GEN_35) : $signed(_GEN_1085); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1169 = 4'h6 == state ? $signed(_GEN_36) : $signed(_GEN_1086); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1170 = 4'h6 == state ? $signed(_GEN_37) : $signed(_GEN_1087); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1171 = 4'h6 == state ? $signed(_GEN_38) : $signed(_GEN_1088); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1172 = 4'h6 == state ? $signed(_GEN_39) : $signed(_GEN_1089); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1173 = 4'h6 == state ? $signed(_GEN_40) : $signed(_GEN_1090); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1174 = 4'h6 == state ? $signed(_GEN_41) : $signed(_GEN_1091); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1175 = 4'h6 == state ? $signed(_GEN_42) : $signed(_GEN_1092); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1176 = 4'h6 == state ? $signed(_GEN_43) : $signed(_GEN_1093); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1177 = 4'h6 == state ? $signed(_GEN_44) : $signed(_GEN_1094); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1178 = 4'h6 == state ? $signed(_GEN_45) : $signed(_GEN_1095); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1179 = 4'h6 == state ? $signed(_GEN_46) : $signed(_GEN_1096); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1180 = 4'h6 == state ? $signed(_GEN_47) : $signed(_GEN_1097); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1181 = 4'h6 == state ? $signed(_GEN_48) : $signed(_GEN_1098); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1182 = 4'h6 == state ? $signed(_GEN_49) : $signed(_GEN_1099); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1183 = 4'h6 == state ? $signed(_GEN_50) : $signed(_GEN_1100); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1184 = 4'h6 == state ? $signed(_GEN_51) : $signed(_GEN_1101); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1185 = 4'h6 == state ? $signed(_GEN_52) : $signed(_GEN_1102); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1186 = 4'h6 == state ? $signed(_GEN_53) : $signed(_GEN_1103); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1187 = 4'h6 == state ? $signed(_GEN_54) : $signed(_GEN_1104); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1188 = 4'h6 == state ? $signed(_GEN_55) : $signed(_GEN_1105); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1189 = 4'h6 == state ? $signed(_GEN_56) : $signed(_GEN_1106); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1190 = 4'h6 == state ? $signed(_GEN_57) : $signed(_GEN_1107); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1191 = 4'h6 == state ? $signed(_GEN_58) : $signed(_GEN_1108); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1192 = 4'h6 == state ? $signed(_GEN_59) : $signed(_GEN_1109); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1193 = 4'h6 == state ? $signed(_GEN_60) : $signed(_GEN_1110); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1194 = 4'h6 == state ? $signed(_GEN_61) : $signed(_GEN_1111); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1195 = 4'h6 == state ? $signed(_GEN_62) : $signed(_GEN_1112); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1196 = 4'h6 == state ? $signed(_GEN_63) : $signed(_GEN_1113); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1197 = 4'h6 == state ? $signed(_GEN_64) : $signed(_GEN_1114); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1198 = 4'h6 == state ? $signed(_GEN_65) : $signed(_GEN_1115); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1199 = 4'h6 == state ? $signed(_GEN_66) : $signed(_GEN_1116); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1200 = 4'h6 == state ? $signed(_GEN_67) : $signed(_GEN_1117); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1201 = 4'h6 == state ? $signed(_GEN_68) : $signed(_GEN_1118); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1202 = 4'h6 == state ? $signed(_GEN_69) : $signed(_GEN_1119); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1203 = 4'h6 == state ? $signed(_GEN_70) : $signed(_GEN_1120); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1204 = 4'h6 == state ? $signed(_GEN_71) : $signed(_GEN_1121); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1205 = 4'h6 == state ? $signed(_GEN_72) : $signed(_GEN_1122); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1206 = 4'h6 == state ? $signed(_GEN_73) : $signed(_GEN_1123); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1207 = 4'h6 == state ? $signed(_GEN_74) : $signed(_GEN_1124); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1208 = 4'h6 == state ? $signed(_GEN_75) : $signed(_GEN_1125); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1209 = 4'h6 == state ? $signed(_GEN_76) : $signed(_GEN_1126); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1210 = 4'h6 == state ? $signed(_GEN_77) : $signed(_GEN_1127); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1211 = 4'h6 == state ? $signed(_GEN_78) : $signed(_GEN_1128); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1212 = 4'h6 == state ? $signed(_GEN_79) : $signed(_GEN_1129); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1213 = 4'h6 == state ? $signed(_GEN_80) : $signed(_GEN_1130); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1214 = 4'h6 == state ? $signed(i) : $signed(_GEN_1131); // @[insertSort.scala 22:16 26:19]
  wire [31:0] _GEN_1215 = 4'h5 == state ? $signed(_GEN_241) : $signed(_GEN_1134); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1216 = 4'h5 == state ? $signed(_GEN_242) : $signed(_GEN_1135); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1217 = 4'h5 == state ? $signed(_GEN_243) : $signed(_GEN_1136); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1218 = 4'h5 == state ? $signed(_GEN_244) : $signed(_GEN_1137); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1219 = 4'h5 == state ? $signed(_GEN_245) : $signed(_GEN_1138); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1220 = 4'h5 == state ? $signed(_GEN_246) : $signed(_GEN_1139); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1221 = 4'h5 == state ? $signed(_GEN_247) : $signed(_GEN_1140); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1222 = 4'h5 == state ? $signed(_GEN_248) : $signed(_GEN_1141); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1223 = 4'h5 == state ? $signed(_GEN_249) : $signed(_GEN_1142); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1224 = 4'h5 == state ? $signed(_GEN_250) : $signed(_GEN_1143); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1225 = 4'h5 == state ? $signed(_GEN_251) : $signed(_GEN_1144); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1226 = 4'h5 == state ? $signed(_GEN_252) : $signed(_GEN_1145); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1227 = 4'h5 == state ? $signed(_GEN_253) : $signed(_GEN_1146); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1228 = 4'h5 == state ? $signed(_GEN_254) : $signed(_GEN_1147); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1229 = 4'h5 == state ? $signed(_GEN_255) : $signed(_GEN_1148); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1230 = 4'h5 == state ? $signed(_GEN_256) : $signed(_GEN_1149); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1231 = 4'h5 == state ? $signed(_GEN_257) : $signed(_GEN_1150); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1232 = 4'h5 == state ? $signed(_GEN_258) : $signed(_GEN_1151); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1233 = 4'h5 == state ? $signed(_GEN_259) : $signed(_GEN_1152); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1234 = 4'h5 == state ? $signed(_GEN_260) : $signed(_GEN_1153); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1235 = 4'h5 == state ? $signed(_GEN_261) : $signed(_GEN_1154); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1236 = 4'h5 == state ? $signed(_GEN_262) : $signed(_GEN_1155); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1237 = 4'h5 == state ? $signed(_GEN_263) : $signed(_GEN_1156); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1238 = 4'h5 == state ? $signed(_GEN_264) : $signed(_GEN_1157); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1239 = 4'h5 == state ? $signed(_GEN_265) : $signed(_GEN_1158); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1240 = 4'h5 == state ? $signed(_GEN_266) : $signed(_GEN_1159); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1241 = 4'h5 == state ? $signed(_GEN_267) : $signed(_GEN_1160); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1242 = 4'h5 == state ? $signed(_GEN_268) : $signed(_GEN_1161); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1243 = 4'h5 == state ? $signed(_GEN_269) : $signed(_GEN_1162); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1244 = 4'h5 == state ? $signed(_GEN_270) : $signed(_GEN_1163); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1245 = 4'h5 == state ? $signed(_GEN_271) : $signed(_GEN_1164); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1246 = 4'h5 == state ? $signed(_GEN_272) : $signed(_GEN_1165); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1247 = 4'h5 == state ? $signed(_GEN_273) : $signed(_GEN_1166); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1248 = 4'h5 == state ? $signed(_GEN_274) : $signed(_GEN_1167); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1249 = 4'h5 == state ? $signed(_GEN_275) : $signed(_GEN_1168); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1250 = 4'h5 == state ? $signed(_GEN_276) : $signed(_GEN_1169); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1251 = 4'h5 == state ? $signed(_GEN_277) : $signed(_GEN_1170); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1252 = 4'h5 == state ? $signed(_GEN_278) : $signed(_GEN_1171); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1253 = 4'h5 == state ? $signed(_GEN_279) : $signed(_GEN_1172); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1254 = 4'h5 == state ? $signed(_GEN_280) : $signed(_GEN_1173); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1255 = 4'h5 == state ? $signed(_GEN_281) : $signed(_GEN_1174); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1256 = 4'h5 == state ? $signed(_GEN_282) : $signed(_GEN_1175); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1257 = 4'h5 == state ? $signed(_GEN_283) : $signed(_GEN_1176); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1258 = 4'h5 == state ? $signed(_GEN_284) : $signed(_GEN_1177); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1259 = 4'h5 == state ? $signed(_GEN_285) : $signed(_GEN_1178); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1260 = 4'h5 == state ? $signed(_GEN_286) : $signed(_GEN_1179); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1261 = 4'h5 == state ? $signed(_GEN_287) : $signed(_GEN_1180); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1262 = 4'h5 == state ? $signed(_GEN_288) : $signed(_GEN_1181); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1263 = 4'h5 == state ? $signed(_GEN_289) : $signed(_GEN_1182); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1264 = 4'h5 == state ? $signed(_GEN_290) : $signed(_GEN_1183); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1265 = 4'h5 == state ? $signed(_GEN_291) : $signed(_GEN_1184); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1266 = 4'h5 == state ? $signed(_GEN_292) : $signed(_GEN_1185); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1267 = 4'h5 == state ? $signed(_GEN_293) : $signed(_GEN_1186); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1268 = 4'h5 == state ? $signed(_GEN_294) : $signed(_GEN_1187); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1269 = 4'h5 == state ? $signed(_GEN_295) : $signed(_GEN_1188); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1270 = 4'h5 == state ? $signed(_GEN_296) : $signed(_GEN_1189); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1271 = 4'h5 == state ? $signed(_GEN_297) : $signed(_GEN_1190); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1272 = 4'h5 == state ? $signed(_GEN_298) : $signed(_GEN_1191); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1273 = 4'h5 == state ? $signed(_GEN_299) : $signed(_GEN_1192); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1274 = 4'h5 == state ? $signed(_GEN_300) : $signed(_GEN_1193); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1275 = 4'h5 == state ? $signed(_GEN_301) : $signed(_GEN_1194); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1276 = 4'h5 == state ? $signed(_GEN_302) : $signed(_GEN_1195); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1277 = 4'h5 == state ? $signed(_GEN_303) : $signed(_GEN_1196); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1278 = 4'h5 == state ? $signed(_GEN_304) : $signed(_GEN_1197); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1279 = 4'h5 == state ? $signed(_GEN_305) : $signed(_GEN_1198); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1280 = 4'h5 == state ? $signed(_GEN_306) : $signed(_GEN_1199); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1281 = 4'h5 == state ? $signed(_GEN_307) : $signed(_GEN_1200); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1282 = 4'h5 == state ? $signed(_GEN_308) : $signed(_GEN_1201); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1283 = 4'h5 == state ? $signed(_GEN_309) : $signed(_GEN_1202); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1284 = 4'h5 == state ? $signed(_GEN_310) : $signed(_GEN_1203); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1285 = 4'h5 == state ? $signed(_GEN_311) : $signed(_GEN_1204); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1286 = 4'h5 == state ? $signed(_GEN_312) : $signed(_GEN_1205); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1287 = 4'h5 == state ? $signed(_GEN_313) : $signed(_GEN_1206); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1288 = 4'h5 == state ? $signed(_GEN_314) : $signed(_GEN_1207); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1289 = 4'h5 == state ? $signed(_GEN_315) : $signed(_GEN_1208); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1290 = 4'h5 == state ? $signed(_GEN_316) : $signed(_GEN_1209); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1291 = 4'h5 == state ? $signed(_GEN_317) : $signed(_GEN_1210); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1292 = 4'h5 == state ? $signed(_GEN_318) : $signed(_GEN_1211); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1293 = 4'h5 == state ? $signed(_GEN_319) : $signed(_GEN_1212); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1294 = 4'h5 == state ? $signed(_GEN_320) : $signed(_GEN_1213); // @[insertSort.scala 26:19]
  wire [3:0] _GEN_1295 = 4'h5 == state ? 4'h6 : _GEN_1133; // @[insertSort.scala 26:19 50:19]
  wire [31:0] _GEN_1296 = 4'h5 == state ? $signed(j) : $signed(_GEN_1132); // @[insertSort.scala 24:16 26:19]
  wire [31:0] _GEN_1297 = 4'h5 == state ? $signed(i) : $signed(_GEN_1214); // @[insertSort.scala 22:16 26:19]
  wire [3:0] _GEN_1298 = 4'h4 == state ? {{1'd0}, _state_T_8} : _GEN_1295; // @[insertSort.scala 26:19 46:19]
  wire [31:0] _GEN_1299 = 4'h4 == state ? $signed(_GEN_1) : $signed(_GEN_1215); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1300 = 4'h4 == state ? $signed(_GEN_2) : $signed(_GEN_1216); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1301 = 4'h4 == state ? $signed(_GEN_3) : $signed(_GEN_1217); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1302 = 4'h4 == state ? $signed(_GEN_4) : $signed(_GEN_1218); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1303 = 4'h4 == state ? $signed(_GEN_5) : $signed(_GEN_1219); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1304 = 4'h4 == state ? $signed(_GEN_6) : $signed(_GEN_1220); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1305 = 4'h4 == state ? $signed(_GEN_7) : $signed(_GEN_1221); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1306 = 4'h4 == state ? $signed(_GEN_8) : $signed(_GEN_1222); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1307 = 4'h4 == state ? $signed(_GEN_9) : $signed(_GEN_1223); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1308 = 4'h4 == state ? $signed(_GEN_10) : $signed(_GEN_1224); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1309 = 4'h4 == state ? $signed(_GEN_11) : $signed(_GEN_1225); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1310 = 4'h4 == state ? $signed(_GEN_12) : $signed(_GEN_1226); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1311 = 4'h4 == state ? $signed(_GEN_13) : $signed(_GEN_1227); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1312 = 4'h4 == state ? $signed(_GEN_14) : $signed(_GEN_1228); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1313 = 4'h4 == state ? $signed(_GEN_15) : $signed(_GEN_1229); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1314 = 4'h4 == state ? $signed(_GEN_16) : $signed(_GEN_1230); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1315 = 4'h4 == state ? $signed(_GEN_17) : $signed(_GEN_1231); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1316 = 4'h4 == state ? $signed(_GEN_18) : $signed(_GEN_1232); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1317 = 4'h4 == state ? $signed(_GEN_19) : $signed(_GEN_1233); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1318 = 4'h4 == state ? $signed(_GEN_20) : $signed(_GEN_1234); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1319 = 4'h4 == state ? $signed(_GEN_21) : $signed(_GEN_1235); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1320 = 4'h4 == state ? $signed(_GEN_22) : $signed(_GEN_1236); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1321 = 4'h4 == state ? $signed(_GEN_23) : $signed(_GEN_1237); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1322 = 4'h4 == state ? $signed(_GEN_24) : $signed(_GEN_1238); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1323 = 4'h4 == state ? $signed(_GEN_25) : $signed(_GEN_1239); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1324 = 4'h4 == state ? $signed(_GEN_26) : $signed(_GEN_1240); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1325 = 4'h4 == state ? $signed(_GEN_27) : $signed(_GEN_1241); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1326 = 4'h4 == state ? $signed(_GEN_28) : $signed(_GEN_1242); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1327 = 4'h4 == state ? $signed(_GEN_29) : $signed(_GEN_1243); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1328 = 4'h4 == state ? $signed(_GEN_30) : $signed(_GEN_1244); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1329 = 4'h4 == state ? $signed(_GEN_31) : $signed(_GEN_1245); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1330 = 4'h4 == state ? $signed(_GEN_32) : $signed(_GEN_1246); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1331 = 4'h4 == state ? $signed(_GEN_33) : $signed(_GEN_1247); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1332 = 4'h4 == state ? $signed(_GEN_34) : $signed(_GEN_1248); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1333 = 4'h4 == state ? $signed(_GEN_35) : $signed(_GEN_1249); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1334 = 4'h4 == state ? $signed(_GEN_36) : $signed(_GEN_1250); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1335 = 4'h4 == state ? $signed(_GEN_37) : $signed(_GEN_1251); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1336 = 4'h4 == state ? $signed(_GEN_38) : $signed(_GEN_1252); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1337 = 4'h4 == state ? $signed(_GEN_39) : $signed(_GEN_1253); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1338 = 4'h4 == state ? $signed(_GEN_40) : $signed(_GEN_1254); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1339 = 4'h4 == state ? $signed(_GEN_41) : $signed(_GEN_1255); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1340 = 4'h4 == state ? $signed(_GEN_42) : $signed(_GEN_1256); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1341 = 4'h4 == state ? $signed(_GEN_43) : $signed(_GEN_1257); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1342 = 4'h4 == state ? $signed(_GEN_44) : $signed(_GEN_1258); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1343 = 4'h4 == state ? $signed(_GEN_45) : $signed(_GEN_1259); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1344 = 4'h4 == state ? $signed(_GEN_46) : $signed(_GEN_1260); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1345 = 4'h4 == state ? $signed(_GEN_47) : $signed(_GEN_1261); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1346 = 4'h4 == state ? $signed(_GEN_48) : $signed(_GEN_1262); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1347 = 4'h4 == state ? $signed(_GEN_49) : $signed(_GEN_1263); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1348 = 4'h4 == state ? $signed(_GEN_50) : $signed(_GEN_1264); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1349 = 4'h4 == state ? $signed(_GEN_51) : $signed(_GEN_1265); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1350 = 4'h4 == state ? $signed(_GEN_52) : $signed(_GEN_1266); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1351 = 4'h4 == state ? $signed(_GEN_53) : $signed(_GEN_1267); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1352 = 4'h4 == state ? $signed(_GEN_54) : $signed(_GEN_1268); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1353 = 4'h4 == state ? $signed(_GEN_55) : $signed(_GEN_1269); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1354 = 4'h4 == state ? $signed(_GEN_56) : $signed(_GEN_1270); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1355 = 4'h4 == state ? $signed(_GEN_57) : $signed(_GEN_1271); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1356 = 4'h4 == state ? $signed(_GEN_58) : $signed(_GEN_1272); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1357 = 4'h4 == state ? $signed(_GEN_59) : $signed(_GEN_1273); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1358 = 4'h4 == state ? $signed(_GEN_60) : $signed(_GEN_1274); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1359 = 4'h4 == state ? $signed(_GEN_61) : $signed(_GEN_1275); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1360 = 4'h4 == state ? $signed(_GEN_62) : $signed(_GEN_1276); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1361 = 4'h4 == state ? $signed(_GEN_63) : $signed(_GEN_1277); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1362 = 4'h4 == state ? $signed(_GEN_64) : $signed(_GEN_1278); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1363 = 4'h4 == state ? $signed(_GEN_65) : $signed(_GEN_1279); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1364 = 4'h4 == state ? $signed(_GEN_66) : $signed(_GEN_1280); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1365 = 4'h4 == state ? $signed(_GEN_67) : $signed(_GEN_1281); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1366 = 4'h4 == state ? $signed(_GEN_68) : $signed(_GEN_1282); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1367 = 4'h4 == state ? $signed(_GEN_69) : $signed(_GEN_1283); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1368 = 4'h4 == state ? $signed(_GEN_70) : $signed(_GEN_1284); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1369 = 4'h4 == state ? $signed(_GEN_71) : $signed(_GEN_1285); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1370 = 4'h4 == state ? $signed(_GEN_72) : $signed(_GEN_1286); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1371 = 4'h4 == state ? $signed(_GEN_73) : $signed(_GEN_1287); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1372 = 4'h4 == state ? $signed(_GEN_74) : $signed(_GEN_1288); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1373 = 4'h4 == state ? $signed(_GEN_75) : $signed(_GEN_1289); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1374 = 4'h4 == state ? $signed(_GEN_76) : $signed(_GEN_1290); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1375 = 4'h4 == state ? $signed(_GEN_77) : $signed(_GEN_1291); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1376 = 4'h4 == state ? $signed(_GEN_78) : $signed(_GEN_1292); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1377 = 4'h4 == state ? $signed(_GEN_79) : $signed(_GEN_1293); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1378 = 4'h4 == state ? $signed(_GEN_80) : $signed(_GEN_1294); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1379 = 4'h4 == state ? $signed(j) : $signed(_GEN_1296); // @[insertSort.scala 24:16 26:19]
  wire [31:0] _GEN_1380 = 4'h4 == state ? $signed(i) : $signed(_GEN_1297); // @[insertSort.scala 22:16 26:19]
  wire [31:0] _GEN_1381 = 4'h3 == state ? $signed(_j_T_2) : $signed(_GEN_1379); // @[insertSort.scala 26:19 42:15]
  wire [3:0] _GEN_1382 = 4'h3 == state ? 4'h4 : _GEN_1298; // @[insertSort.scala 26:19 43:19]
  wire [31:0] _GEN_1383 = 4'h3 == state ? $signed(_GEN_1) : $signed(_GEN_1299); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1384 = 4'h3 == state ? $signed(_GEN_2) : $signed(_GEN_1300); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1385 = 4'h3 == state ? $signed(_GEN_3) : $signed(_GEN_1301); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1386 = 4'h3 == state ? $signed(_GEN_4) : $signed(_GEN_1302); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1387 = 4'h3 == state ? $signed(_GEN_5) : $signed(_GEN_1303); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1388 = 4'h3 == state ? $signed(_GEN_6) : $signed(_GEN_1304); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1389 = 4'h3 == state ? $signed(_GEN_7) : $signed(_GEN_1305); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1390 = 4'h3 == state ? $signed(_GEN_8) : $signed(_GEN_1306); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1391 = 4'h3 == state ? $signed(_GEN_9) : $signed(_GEN_1307); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1392 = 4'h3 == state ? $signed(_GEN_10) : $signed(_GEN_1308); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1393 = 4'h3 == state ? $signed(_GEN_11) : $signed(_GEN_1309); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1394 = 4'h3 == state ? $signed(_GEN_12) : $signed(_GEN_1310); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1395 = 4'h3 == state ? $signed(_GEN_13) : $signed(_GEN_1311); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1396 = 4'h3 == state ? $signed(_GEN_14) : $signed(_GEN_1312); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1397 = 4'h3 == state ? $signed(_GEN_15) : $signed(_GEN_1313); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1398 = 4'h3 == state ? $signed(_GEN_16) : $signed(_GEN_1314); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1399 = 4'h3 == state ? $signed(_GEN_17) : $signed(_GEN_1315); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1400 = 4'h3 == state ? $signed(_GEN_18) : $signed(_GEN_1316); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1401 = 4'h3 == state ? $signed(_GEN_19) : $signed(_GEN_1317); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1402 = 4'h3 == state ? $signed(_GEN_20) : $signed(_GEN_1318); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1403 = 4'h3 == state ? $signed(_GEN_21) : $signed(_GEN_1319); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1404 = 4'h3 == state ? $signed(_GEN_22) : $signed(_GEN_1320); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1405 = 4'h3 == state ? $signed(_GEN_23) : $signed(_GEN_1321); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1406 = 4'h3 == state ? $signed(_GEN_24) : $signed(_GEN_1322); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1407 = 4'h3 == state ? $signed(_GEN_25) : $signed(_GEN_1323); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1408 = 4'h3 == state ? $signed(_GEN_26) : $signed(_GEN_1324); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1409 = 4'h3 == state ? $signed(_GEN_27) : $signed(_GEN_1325); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1410 = 4'h3 == state ? $signed(_GEN_28) : $signed(_GEN_1326); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1411 = 4'h3 == state ? $signed(_GEN_29) : $signed(_GEN_1327); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1412 = 4'h3 == state ? $signed(_GEN_30) : $signed(_GEN_1328); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1413 = 4'h3 == state ? $signed(_GEN_31) : $signed(_GEN_1329); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1414 = 4'h3 == state ? $signed(_GEN_32) : $signed(_GEN_1330); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1415 = 4'h3 == state ? $signed(_GEN_33) : $signed(_GEN_1331); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1416 = 4'h3 == state ? $signed(_GEN_34) : $signed(_GEN_1332); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1417 = 4'h3 == state ? $signed(_GEN_35) : $signed(_GEN_1333); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1418 = 4'h3 == state ? $signed(_GEN_36) : $signed(_GEN_1334); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1419 = 4'h3 == state ? $signed(_GEN_37) : $signed(_GEN_1335); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1420 = 4'h3 == state ? $signed(_GEN_38) : $signed(_GEN_1336); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1421 = 4'h3 == state ? $signed(_GEN_39) : $signed(_GEN_1337); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1422 = 4'h3 == state ? $signed(_GEN_40) : $signed(_GEN_1338); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1423 = 4'h3 == state ? $signed(_GEN_41) : $signed(_GEN_1339); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1424 = 4'h3 == state ? $signed(_GEN_42) : $signed(_GEN_1340); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1425 = 4'h3 == state ? $signed(_GEN_43) : $signed(_GEN_1341); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1426 = 4'h3 == state ? $signed(_GEN_44) : $signed(_GEN_1342); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1427 = 4'h3 == state ? $signed(_GEN_45) : $signed(_GEN_1343); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1428 = 4'h3 == state ? $signed(_GEN_46) : $signed(_GEN_1344); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1429 = 4'h3 == state ? $signed(_GEN_47) : $signed(_GEN_1345); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1430 = 4'h3 == state ? $signed(_GEN_48) : $signed(_GEN_1346); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1431 = 4'h3 == state ? $signed(_GEN_49) : $signed(_GEN_1347); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1432 = 4'h3 == state ? $signed(_GEN_50) : $signed(_GEN_1348); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1433 = 4'h3 == state ? $signed(_GEN_51) : $signed(_GEN_1349); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1434 = 4'h3 == state ? $signed(_GEN_52) : $signed(_GEN_1350); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1435 = 4'h3 == state ? $signed(_GEN_53) : $signed(_GEN_1351); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1436 = 4'h3 == state ? $signed(_GEN_54) : $signed(_GEN_1352); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1437 = 4'h3 == state ? $signed(_GEN_55) : $signed(_GEN_1353); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1438 = 4'h3 == state ? $signed(_GEN_56) : $signed(_GEN_1354); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1439 = 4'h3 == state ? $signed(_GEN_57) : $signed(_GEN_1355); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1440 = 4'h3 == state ? $signed(_GEN_58) : $signed(_GEN_1356); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1441 = 4'h3 == state ? $signed(_GEN_59) : $signed(_GEN_1357); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1442 = 4'h3 == state ? $signed(_GEN_60) : $signed(_GEN_1358); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1443 = 4'h3 == state ? $signed(_GEN_61) : $signed(_GEN_1359); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1444 = 4'h3 == state ? $signed(_GEN_62) : $signed(_GEN_1360); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1445 = 4'h3 == state ? $signed(_GEN_63) : $signed(_GEN_1361); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1446 = 4'h3 == state ? $signed(_GEN_64) : $signed(_GEN_1362); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1447 = 4'h3 == state ? $signed(_GEN_65) : $signed(_GEN_1363); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1448 = 4'h3 == state ? $signed(_GEN_66) : $signed(_GEN_1364); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1449 = 4'h3 == state ? $signed(_GEN_67) : $signed(_GEN_1365); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1450 = 4'h3 == state ? $signed(_GEN_68) : $signed(_GEN_1366); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1451 = 4'h3 == state ? $signed(_GEN_69) : $signed(_GEN_1367); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1452 = 4'h3 == state ? $signed(_GEN_70) : $signed(_GEN_1368); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1453 = 4'h3 == state ? $signed(_GEN_71) : $signed(_GEN_1369); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1454 = 4'h3 == state ? $signed(_GEN_72) : $signed(_GEN_1370); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1455 = 4'h3 == state ? $signed(_GEN_73) : $signed(_GEN_1371); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1456 = 4'h3 == state ? $signed(_GEN_74) : $signed(_GEN_1372); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1457 = 4'h3 == state ? $signed(_GEN_75) : $signed(_GEN_1373); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1458 = 4'h3 == state ? $signed(_GEN_76) : $signed(_GEN_1374); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1459 = 4'h3 == state ? $signed(_GEN_77) : $signed(_GEN_1375); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1460 = 4'h3 == state ? $signed(_GEN_78) : $signed(_GEN_1376); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1461 = 4'h3 == state ? $signed(_GEN_79) : $signed(_GEN_1377); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1462 = 4'h3 == state ? $signed(_GEN_80) : $signed(_GEN_1378); // @[insertSort.scala 26:19]
  wire [31:0] _GEN_1463 = 4'h3 == state ? $signed(i) : $signed(_GEN_1380); // @[insertSort.scala 22:16 26:19]
  wire [3:0] _GEN_1465 = 4'h2 == state ? 4'h3 : _GEN_1382; // @[insertSort.scala 26:19 39:19]
  assign io_array_out_0 = array_0; // @[insertSort.scala 21:18]
  assign io_array_out_1 = array_1; // @[insertSort.scala 21:18]
  assign io_array_out_2 = array_2; // @[insertSort.scala 21:18]
  assign io_array_out_3 = array_3; // @[insertSort.scala 21:18]
  assign io_array_out_4 = array_4; // @[insertSort.scala 21:18]
  assign io_array_out_5 = array_5; // @[insertSort.scala 21:18]
  assign io_array_out_6 = array_6; // @[insertSort.scala 21:18]
  assign io_array_out_7 = array_7; // @[insertSort.scala 21:18]
  assign io_array_out_8 = array_8; // @[insertSort.scala 21:18]
  assign io_array_out_9 = array_9; // @[insertSort.scala 21:18]
  assign io_array_out_10 = array_10; // @[insertSort.scala 21:18]
  assign io_array_out_11 = array_11; // @[insertSort.scala 21:18]
  assign io_array_out_12 = array_12; // @[insertSort.scala 21:18]
  assign io_array_out_13 = array_13; // @[insertSort.scala 21:18]
  assign io_array_out_14 = array_14; // @[insertSort.scala 21:18]
  assign io_array_out_15 = array_15; // @[insertSort.scala 21:18]
  assign io_array_out_16 = array_16; // @[insertSort.scala 21:18]
  assign io_array_out_17 = array_17; // @[insertSort.scala 21:18]
  assign io_array_out_18 = array_18; // @[insertSort.scala 21:18]
  assign io_array_out_19 = array_19; // @[insertSort.scala 21:18]
  assign io_ready = state == 4'hc; // @[insertSort.scala 80:23]
  always @(posedge clock) begin
    if (reset) begin // @[insertSort.scala 13:24]
      state <= 4'hf; // @[insertSort.scala 13:24]
    end else if (4'hf == state) begin // @[insertSort.scala 26:19]
      if (io_valid) begin // @[insertSort.scala 28:25]
        state <= 4'h0;
      end
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      state <= 4'h1; // @[insertSort.scala 32:19]
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      state <= _state_T_2; // @[insertSort.scala 35:19]
    end else begin
      state <= _GEN_1465;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_0 <= _GEN_1;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_0 <= _GEN_1;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_0 <= _GEN_1;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_0 <= _GEN_1;
    end else begin
      array_0 <= _GEN_1383;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_1 <= _GEN_2;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_1 <= _GEN_2;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_1 <= _GEN_2;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_1 <= _GEN_2;
    end else begin
      array_1 <= _GEN_1384;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_2 <= _GEN_3;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_2 <= _GEN_3;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_2 <= _GEN_3;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_2 <= _GEN_3;
    end else begin
      array_2 <= _GEN_1385;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_3 <= _GEN_4;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_3 <= _GEN_4;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_3 <= _GEN_4;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_3 <= _GEN_4;
    end else begin
      array_3 <= _GEN_1386;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_4 <= _GEN_5;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_4 <= _GEN_5;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_4 <= _GEN_5;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_4 <= _GEN_5;
    end else begin
      array_4 <= _GEN_1387;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_5 <= _GEN_6;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_5 <= _GEN_6;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_5 <= _GEN_6;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_5 <= _GEN_6;
    end else begin
      array_5 <= _GEN_1388;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_6 <= _GEN_7;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_6 <= _GEN_7;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_6 <= _GEN_7;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_6 <= _GEN_7;
    end else begin
      array_6 <= _GEN_1389;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_7 <= _GEN_8;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_7 <= _GEN_8;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_7 <= _GEN_8;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_7 <= _GEN_8;
    end else begin
      array_7 <= _GEN_1390;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_8 <= _GEN_9;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_8 <= _GEN_9;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_8 <= _GEN_9;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_8 <= _GEN_9;
    end else begin
      array_8 <= _GEN_1391;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_9 <= _GEN_10;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_9 <= _GEN_10;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_9 <= _GEN_10;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_9 <= _GEN_10;
    end else begin
      array_9 <= _GEN_1392;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_10 <= _GEN_11;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_10 <= _GEN_11;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_10 <= _GEN_11;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_10 <= _GEN_11;
    end else begin
      array_10 <= _GEN_1393;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_11 <= _GEN_12;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_11 <= _GEN_12;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_11 <= _GEN_12;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_11 <= _GEN_12;
    end else begin
      array_11 <= _GEN_1394;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_12 <= _GEN_13;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_12 <= _GEN_13;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_12 <= _GEN_13;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_12 <= _GEN_13;
    end else begin
      array_12 <= _GEN_1395;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_13 <= _GEN_14;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_13 <= _GEN_14;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_13 <= _GEN_14;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_13 <= _GEN_14;
    end else begin
      array_13 <= _GEN_1396;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_14 <= _GEN_15;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_14 <= _GEN_15;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_14 <= _GEN_15;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_14 <= _GEN_15;
    end else begin
      array_14 <= _GEN_1397;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_15 <= _GEN_16;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_15 <= _GEN_16;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_15 <= _GEN_16;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_15 <= _GEN_16;
    end else begin
      array_15 <= _GEN_1398;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_16 <= _GEN_17;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_16 <= _GEN_17;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_16 <= _GEN_17;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_16 <= _GEN_17;
    end else begin
      array_16 <= _GEN_1399;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_17 <= _GEN_18;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_17 <= _GEN_18;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_17 <= _GEN_18;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_17 <= _GEN_18;
    end else begin
      array_17 <= _GEN_1400;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_18 <= _GEN_19;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_18 <= _GEN_19;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_18 <= _GEN_19;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_18 <= _GEN_19;
    end else begin
      array_18 <= _GEN_1401;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_19 <= _GEN_20;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_19 <= _GEN_20;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_19 <= _GEN_20;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_19 <= _GEN_20;
    end else begin
      array_19 <= _GEN_1402;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_20 <= _GEN_21;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_20 <= _GEN_21;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_20 <= _GEN_21;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_20 <= _GEN_21;
    end else begin
      array_20 <= _GEN_1403;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_21 <= _GEN_22;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_21 <= _GEN_22;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_21 <= _GEN_22;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_21 <= _GEN_22;
    end else begin
      array_21 <= _GEN_1404;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_22 <= _GEN_23;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_22 <= _GEN_23;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_22 <= _GEN_23;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_22 <= _GEN_23;
    end else begin
      array_22 <= _GEN_1405;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_23 <= _GEN_24;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_23 <= _GEN_24;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_23 <= _GEN_24;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_23 <= _GEN_24;
    end else begin
      array_23 <= _GEN_1406;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_24 <= _GEN_25;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_24 <= _GEN_25;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_24 <= _GEN_25;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_24 <= _GEN_25;
    end else begin
      array_24 <= _GEN_1407;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_25 <= _GEN_26;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_25 <= _GEN_26;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_25 <= _GEN_26;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_25 <= _GEN_26;
    end else begin
      array_25 <= _GEN_1408;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_26 <= _GEN_27;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_26 <= _GEN_27;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_26 <= _GEN_27;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_26 <= _GEN_27;
    end else begin
      array_26 <= _GEN_1409;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_27 <= _GEN_28;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_27 <= _GEN_28;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_27 <= _GEN_28;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_27 <= _GEN_28;
    end else begin
      array_27 <= _GEN_1410;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_28 <= _GEN_29;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_28 <= _GEN_29;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_28 <= _GEN_29;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_28 <= _GEN_29;
    end else begin
      array_28 <= _GEN_1411;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_29 <= _GEN_30;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_29 <= _GEN_30;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_29 <= _GEN_30;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_29 <= _GEN_30;
    end else begin
      array_29 <= _GEN_1412;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_30 <= _GEN_31;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_30 <= _GEN_31;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_30 <= _GEN_31;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_30 <= _GEN_31;
    end else begin
      array_30 <= _GEN_1413;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_31 <= _GEN_32;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_31 <= _GEN_32;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_31 <= _GEN_32;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_31 <= _GEN_32;
    end else begin
      array_31 <= _GEN_1414;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_32 <= _GEN_33;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_32 <= _GEN_33;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_32 <= _GEN_33;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_32 <= _GEN_33;
    end else begin
      array_32 <= _GEN_1415;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_33 <= _GEN_34;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_33 <= _GEN_34;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_33 <= _GEN_34;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_33 <= _GEN_34;
    end else begin
      array_33 <= _GEN_1416;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_34 <= _GEN_35;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_34 <= _GEN_35;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_34 <= _GEN_35;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_34 <= _GEN_35;
    end else begin
      array_34 <= _GEN_1417;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_35 <= _GEN_36;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_35 <= _GEN_36;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_35 <= _GEN_36;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_35 <= _GEN_36;
    end else begin
      array_35 <= _GEN_1418;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_36 <= _GEN_37;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_36 <= _GEN_37;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_36 <= _GEN_37;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_36 <= _GEN_37;
    end else begin
      array_36 <= _GEN_1419;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_37 <= _GEN_38;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_37 <= _GEN_38;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_37 <= _GEN_38;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_37 <= _GEN_38;
    end else begin
      array_37 <= _GEN_1420;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_38 <= _GEN_39;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_38 <= _GEN_39;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_38 <= _GEN_39;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_38 <= _GEN_39;
    end else begin
      array_38 <= _GEN_1421;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_39 <= _GEN_40;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_39 <= _GEN_40;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_39 <= _GEN_40;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_39 <= _GEN_40;
    end else begin
      array_39 <= _GEN_1422;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_40 <= _GEN_41;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_40 <= _GEN_41;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_40 <= _GEN_41;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_40 <= _GEN_41;
    end else begin
      array_40 <= _GEN_1423;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_41 <= _GEN_42;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_41 <= _GEN_42;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_41 <= _GEN_42;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_41 <= _GEN_42;
    end else begin
      array_41 <= _GEN_1424;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_42 <= _GEN_43;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_42 <= _GEN_43;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_42 <= _GEN_43;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_42 <= _GEN_43;
    end else begin
      array_42 <= _GEN_1425;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_43 <= _GEN_44;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_43 <= _GEN_44;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_43 <= _GEN_44;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_43 <= _GEN_44;
    end else begin
      array_43 <= _GEN_1426;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_44 <= _GEN_45;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_44 <= _GEN_45;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_44 <= _GEN_45;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_44 <= _GEN_45;
    end else begin
      array_44 <= _GEN_1427;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_45 <= _GEN_46;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_45 <= _GEN_46;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_45 <= _GEN_46;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_45 <= _GEN_46;
    end else begin
      array_45 <= _GEN_1428;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_46 <= _GEN_47;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_46 <= _GEN_47;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_46 <= _GEN_47;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_46 <= _GEN_47;
    end else begin
      array_46 <= _GEN_1429;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_47 <= _GEN_48;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_47 <= _GEN_48;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_47 <= _GEN_48;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_47 <= _GEN_48;
    end else begin
      array_47 <= _GEN_1430;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_48 <= _GEN_49;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_48 <= _GEN_49;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_48 <= _GEN_49;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_48 <= _GEN_49;
    end else begin
      array_48 <= _GEN_1431;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_49 <= _GEN_50;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_49 <= _GEN_50;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_49 <= _GEN_50;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_49 <= _GEN_50;
    end else begin
      array_49 <= _GEN_1432;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_50 <= _GEN_51;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_50 <= _GEN_51;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_50 <= _GEN_51;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_50 <= _GEN_51;
    end else begin
      array_50 <= _GEN_1433;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_51 <= _GEN_52;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_51 <= _GEN_52;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_51 <= _GEN_52;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_51 <= _GEN_52;
    end else begin
      array_51 <= _GEN_1434;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_52 <= _GEN_53;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_52 <= _GEN_53;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_52 <= _GEN_53;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_52 <= _GEN_53;
    end else begin
      array_52 <= _GEN_1435;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_53 <= _GEN_54;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_53 <= _GEN_54;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_53 <= _GEN_54;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_53 <= _GEN_54;
    end else begin
      array_53 <= _GEN_1436;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_54 <= _GEN_55;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_54 <= _GEN_55;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_54 <= _GEN_55;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_54 <= _GEN_55;
    end else begin
      array_54 <= _GEN_1437;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_55 <= _GEN_56;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_55 <= _GEN_56;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_55 <= _GEN_56;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_55 <= _GEN_56;
    end else begin
      array_55 <= _GEN_1438;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_56 <= _GEN_57;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_56 <= _GEN_57;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_56 <= _GEN_57;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_56 <= _GEN_57;
    end else begin
      array_56 <= _GEN_1439;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_57 <= _GEN_58;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_57 <= _GEN_58;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_57 <= _GEN_58;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_57 <= _GEN_58;
    end else begin
      array_57 <= _GEN_1440;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_58 <= _GEN_59;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_58 <= _GEN_59;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_58 <= _GEN_59;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_58 <= _GEN_59;
    end else begin
      array_58 <= _GEN_1441;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_59 <= _GEN_60;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_59 <= _GEN_60;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_59 <= _GEN_60;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_59 <= _GEN_60;
    end else begin
      array_59 <= _GEN_1442;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_60 <= _GEN_61;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_60 <= _GEN_61;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_60 <= _GEN_61;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_60 <= _GEN_61;
    end else begin
      array_60 <= _GEN_1443;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_61 <= _GEN_62;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_61 <= _GEN_62;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_61 <= _GEN_62;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_61 <= _GEN_62;
    end else begin
      array_61 <= _GEN_1444;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_62 <= _GEN_63;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_62 <= _GEN_63;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_62 <= _GEN_63;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_62 <= _GEN_63;
    end else begin
      array_62 <= _GEN_1445;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_63 <= _GEN_64;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_63 <= _GEN_64;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_63 <= _GEN_64;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_63 <= _GEN_64;
    end else begin
      array_63 <= _GEN_1446;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_64 <= _GEN_65;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_64 <= _GEN_65;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_64 <= _GEN_65;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_64 <= _GEN_65;
    end else begin
      array_64 <= _GEN_1447;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_65 <= _GEN_66;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_65 <= _GEN_66;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_65 <= _GEN_66;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_65 <= _GEN_66;
    end else begin
      array_65 <= _GEN_1448;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_66 <= _GEN_67;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_66 <= _GEN_67;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_66 <= _GEN_67;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_66 <= _GEN_67;
    end else begin
      array_66 <= _GEN_1449;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_67 <= _GEN_68;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_67 <= _GEN_68;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_67 <= _GEN_68;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_67 <= _GEN_68;
    end else begin
      array_67 <= _GEN_1450;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_68 <= _GEN_69;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_68 <= _GEN_69;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_68 <= _GEN_69;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_68 <= _GEN_69;
    end else begin
      array_68 <= _GEN_1451;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_69 <= _GEN_70;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_69 <= _GEN_70;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_69 <= _GEN_70;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_69 <= _GEN_70;
    end else begin
      array_69 <= _GEN_1452;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_70 <= _GEN_71;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_70 <= _GEN_71;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_70 <= _GEN_71;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_70 <= _GEN_71;
    end else begin
      array_70 <= _GEN_1453;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_71 <= _GEN_72;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_71 <= _GEN_72;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_71 <= _GEN_72;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_71 <= _GEN_72;
    end else begin
      array_71 <= _GEN_1454;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_72 <= _GEN_73;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_72 <= _GEN_73;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_72 <= _GEN_73;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_72 <= _GEN_73;
    end else begin
      array_72 <= _GEN_1455;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_73 <= _GEN_74;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_73 <= _GEN_74;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_73 <= _GEN_74;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_73 <= _GEN_74;
    end else begin
      array_73 <= _GEN_1456;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_74 <= _GEN_75;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_74 <= _GEN_75;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_74 <= _GEN_75;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_74 <= _GEN_75;
    end else begin
      array_74 <= _GEN_1457;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_75 <= _GEN_76;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_75 <= _GEN_76;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_75 <= _GEN_76;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_75 <= _GEN_76;
    end else begin
      array_75 <= _GEN_1458;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_76 <= _GEN_77;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_76 <= _GEN_77;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_76 <= _GEN_77;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_76 <= _GEN_77;
    end else begin
      array_76 <= _GEN_1459;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_77 <= _GEN_78;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_77 <= _GEN_78;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_77 <= _GEN_78;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_77 <= _GEN_78;
    end else begin
      array_77 <= _GEN_1460;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_78 <= _GEN_79;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_78 <= _GEN_79;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_78 <= _GEN_79;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_78 <= _GEN_79;
    end else begin
      array_78 <= _GEN_1461;
    end
    if (4'hf == state) begin // @[insertSort.scala 26:19]
      array_79 <= _GEN_80;
    end else if (4'h0 == state) begin // @[insertSort.scala 26:19]
      array_79 <= _GEN_80;
    end else if (4'h1 == state) begin // @[insertSort.scala 26:19]
      array_79 <= _GEN_80;
    end else if (4'h2 == state) begin // @[insertSort.scala 26:19]
      array_79 <= _GEN_80;
    end else begin
      array_79 <= _GEN_1462;
    end
    REG <= ~io_valid; // @[insertSort.scala 18:18]
    if (!(4'hf == state)) begin // @[insertSort.scala 26:19]
      if (4'h0 == state) begin // @[insertSort.scala 26:19]
        i <= 32'sh1; // @[insertSort.scala 31:15]
      end else if (!(4'h1 == state)) begin // @[insertSort.scala 26:19]
        if (!(4'h2 == state)) begin // @[insertSort.scala 26:19]
          i <= _GEN_1463;
        end
      end
    end
    if (!(4'hf == state)) begin // @[insertSort.scala 26:19]
      if (!(4'h0 == state)) begin // @[insertSort.scala 26:19]
        if (!(4'h1 == state)) begin // @[insertSort.scala 26:19]
          if (4'h2 == state) begin // @[insertSort.scala 26:19]
            key <= _GEN_160; // @[insertSort.scala 38:17]
          end
        end
      end
    end
    if (!(4'hf == state)) begin // @[insertSort.scala 26:19]
      if (!(4'h0 == state)) begin // @[insertSort.scala 26:19]
        if (!(4'h1 == state)) begin // @[insertSort.scala 26:19]
          if (!(4'h2 == state)) begin // @[insertSort.scala 26:19]
            j <= _GEN_1381;
          end
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  array_0 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  array_1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  array_2 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  array_3 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  array_4 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  array_5 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  array_6 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  array_7 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  array_8 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  array_9 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  array_10 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  array_11 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  array_12 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  array_13 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  array_14 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  array_15 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  array_16 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  array_17 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  array_18 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  array_19 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  array_20 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  array_21 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  array_22 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  array_23 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  array_24 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  array_25 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  array_26 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  array_27 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  array_28 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  array_29 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  array_30 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  array_31 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  array_32 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  array_33 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  array_34 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  array_35 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  array_36 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  array_37 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  array_38 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  array_39 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  array_40 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  array_41 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  array_42 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  array_43 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  array_44 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  array_45 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  array_46 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  array_47 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  array_48 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  array_49 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  array_50 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  array_51 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  array_52 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  array_53 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  array_54 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  array_55 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  array_56 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  array_57 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  array_58 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  array_59 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  array_60 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  array_61 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  array_62 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  array_63 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  array_64 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  array_65 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  array_66 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  array_67 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  array_68 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  array_69 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  array_70 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  array_71 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  array_72 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  array_73 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  array_74 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  array_75 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  array_76 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  array_77 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  array_78 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  array_79 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  REG = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  i = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  key = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  j = _RAND_84[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXIWrapperChiselInsertSort(
  input         clock,
  input         reset,
  input  [31:0] io_S_AXI_AWADDR,
  input  [2:0]  io_S_AXI_AWPROT,
  input         io_S_AXI_AWVALID,
  output        io_S_AXI_AWREADY,
  input  [31:0] io_S_AXI_WDATA,
  input  [3:0]  io_S_AXI_WSTRB,
  input         io_S_AXI_WVALID,
  output        io_S_AXI_WREADY,
  output [1:0]  io_S_AXI_BRESP,
  output        io_S_AXI_BVALID,
  input         io_S_AXI_BREADY,
  input  [31:0] io_S_AXI_ARADDR,
  input  [2:0]  io_S_AXI_ARPROT,
  input         io_S_AXI_ARVALID,
  output        io_S_AXI_ARREADY,
  output [31:0] io_S_AXI_RDATA,
  output [1:0]  io_S_AXI_RRESP,
  output        io_S_AXI_RVALID,
  input         io_S_AXI_RREADY
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  wire  modInsertSort_clock; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire  modInsertSort_reset; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_0; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_1; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_2; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_3; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_4; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_5; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_6; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_7; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_8; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_9; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_10; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_11; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_12; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_13; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_14; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_15; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_16; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_17; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_18; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_19; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire  modInsertSort_io_valid; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_out_0; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_out_1; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_out_2; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_out_3; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_out_4; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_out_5; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_out_6; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_out_7; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_out_8; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_out_9; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_out_10; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_out_11; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_out_12; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_out_13; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_out_14; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_out_15; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_out_16; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_out_17; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_out_18; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire [31:0] modInsertSort_io_array_out_19; // @[AXIWrapperChiselInsertSort.scala 40:31]
  wire  modInsertSort_io_ready; // @[AXIWrapperChiselInsertSort.scala 40:31]
  reg [31:0] axi_awaddr; // @[AXIWrapperChiselInsertSort.scala 43:26]
  reg [31:0] axi_araddr; // @[AXIWrapperChiselInsertSort.scala 44:26]
  reg  axi_awready; // @[AXIWrapperChiselInsertSort.scala 46:26]
  reg  axi_wready; // @[AXIWrapperChiselInsertSort.scala 47:26]
  reg  axi_bvalid; // @[AXIWrapperChiselInsertSort.scala 49:26]
  reg  axi_arready; // @[AXIWrapperChiselInsertSort.scala 50:26]
  reg [31:0] axi_rdata; // @[AXIWrapperChiselInsertSort.scala 51:26]
  reg  axi_rvalid; // @[AXIWrapperChiselInsertSort.scala 53:26]
  reg [31:0] io_valid_reg; // @[AXIWrapperChiselInsertSort.scala 67:27]
  reg [7:0] io_array_0; // @[AXIWrapperChiselInsertSort.scala 70:27]
  reg [7:0] io_array_1; // @[AXIWrapperChiselInsertSort.scala 70:27]
  reg [7:0] io_array_2; // @[AXIWrapperChiselInsertSort.scala 70:27]
  reg [7:0] io_array_3; // @[AXIWrapperChiselInsertSort.scala 70:27]
  reg [7:0] io_array_4; // @[AXIWrapperChiselInsertSort.scala 70:27]
  reg [7:0] io_array_5; // @[AXIWrapperChiselInsertSort.scala 70:27]
  reg [7:0] io_array_6; // @[AXIWrapperChiselInsertSort.scala 70:27]
  reg [7:0] io_array_7; // @[AXIWrapperChiselInsertSort.scala 70:27]
  reg [7:0] io_array_8; // @[AXIWrapperChiselInsertSort.scala 70:27]
  reg [7:0] io_array_9; // @[AXIWrapperChiselInsertSort.scala 70:27]
  reg [7:0] io_array_10; // @[AXIWrapperChiselInsertSort.scala 70:27]
  reg [7:0] io_array_11; // @[AXIWrapperChiselInsertSort.scala 70:27]
  reg [7:0] io_array_12; // @[AXIWrapperChiselInsertSort.scala 70:27]
  reg [7:0] io_array_13; // @[AXIWrapperChiselInsertSort.scala 70:27]
  reg [7:0] io_array_14; // @[AXIWrapperChiselInsertSort.scala 70:27]
  reg [7:0] io_array_15; // @[AXIWrapperChiselInsertSort.scala 70:27]
  reg [7:0] io_array_16; // @[AXIWrapperChiselInsertSort.scala 70:27]
  reg [7:0] io_array_17; // @[AXIWrapperChiselInsertSort.scala 70:27]
  reg [7:0] io_array_18; // @[AXIWrapperChiselInsertSort.scala 70:27]
  reg [7:0] io_array_19; // @[AXIWrapperChiselInsertSort.scala 70:27]
  reg [31:0] reg_data_out; // @[AXIWrapperChiselInsertSort.scala 74:27]
  reg  aw_en; // @[AXIWrapperChiselInsertSort.scala 75:27]
  wire  _T_4 = ~axi_awready & io_S_AXI_AWVALID & io_S_AXI_WVALID & aw_en; // @[AXIWrapperChiselInsertSort.scala 95:66]
  wire  _T_5 = io_S_AXI_BREADY & axi_bvalid; // @[AXIWrapperChiselInsertSort.scala 102:37]
  wire  _GEN_1 = io_S_AXI_BREADY & axi_bvalid | aw_en; // @[AXIWrapperChiselInsertSort.scala 102:52 106:25 75:27]
  wire  _GEN_3 = ~axi_awready & io_S_AXI_AWVALID & io_S_AXI_WVALID & aw_en ? 1'h0 : _GEN_1; // @[AXIWrapperChiselInsertSort.scala 101:25 95:76]
  wire  _T_15 = ~axi_wready & io_S_AXI_WVALID & io_S_AXI_AWVALID & aw_en; // @[AXIWrapperChiselInsertSort.scala 130:65]
  wire  slv_reg_wren = axi_wready & io_S_AXI_WVALID & axi_awready & io_S_AXI_AWVALID; // @[AXIWrapperChiselInsertSort.scala 148:66]
  wire [7:0] _io_array_T_20 = io_S_AXI_WDATA[7:0]; // @[AXIWrapperChiselInsertSort.scala 157:{78,78}]
  wire  _GEN_92 = _T_5 ? 1'h0 : axi_bvalid; // @[AXIWrapperChiselInsertSort.scala 175:49 176:28 49:26]
  wire  _GEN_93 = axi_awready & io_S_AXI_AWVALID & ~axi_bvalid & axi_wready & io_S_AXI_WVALID | _GEN_92; // @[AXIWrapperChiselInsertSort.scala 171:95 172:24]
  wire  _T_30 = ~axi_arready & io_S_AXI_ARVALID; // @[AXIWrapperChiselInsertSort.scala 191:27]
  wire  _T_34 = axi_arready & io_S_AXI_ARVALID & ~axi_rvalid; // @[AXIWrapperChiselInsertSort.scala 212:46]
  wire  _GEN_101 = axi_rvalid & io_S_AXI_RREADY ? 1'h0 : axi_rvalid; // @[AXIWrapperChiselInsertSort.scala 215:52 216:24 53:26]
  wire  _GEN_102 = axi_arready & io_S_AXI_ARVALID & ~axi_rvalid | _GEN_101; // @[AXIWrapperChiselInsertSort.scala 212:62 213:24]
  wire  io_ready = modInsertSort_io_ready; // @[AXIWrapperChiselInsertSort.scala 224:14 69:28]
  wire [7:0] readAddr = axi_araddr[9:2]; // @[AXIWrapperChiselInsertSort.scala 246:30]
  wire [7:0] _GEN_108 = 5'h1 == readAddr[4:0] ? $signed(io_array_1) : $signed(io_array_0); // @[AXIWrapperChiselInsertSort.scala 248:{22,22}]
  wire [7:0] _GEN_109 = 5'h2 == readAddr[4:0] ? $signed(io_array_2) : $signed(_GEN_108); // @[AXIWrapperChiselInsertSort.scala 248:{22,22}]
  wire [7:0] _GEN_110 = 5'h3 == readAddr[4:0] ? $signed(io_array_3) : $signed(_GEN_109); // @[AXIWrapperChiselInsertSort.scala 248:{22,22}]
  wire [7:0] _GEN_111 = 5'h4 == readAddr[4:0] ? $signed(io_array_4) : $signed(_GEN_110); // @[AXIWrapperChiselInsertSort.scala 248:{22,22}]
  wire [7:0] _GEN_112 = 5'h5 == readAddr[4:0] ? $signed(io_array_5) : $signed(_GEN_111); // @[AXIWrapperChiselInsertSort.scala 248:{22,22}]
  wire [7:0] _GEN_113 = 5'h6 == readAddr[4:0] ? $signed(io_array_6) : $signed(_GEN_112); // @[AXIWrapperChiselInsertSort.scala 248:{22,22}]
  wire [7:0] _GEN_114 = 5'h7 == readAddr[4:0] ? $signed(io_array_7) : $signed(_GEN_113); // @[AXIWrapperChiselInsertSort.scala 248:{22,22}]
  wire [7:0] _GEN_115 = 5'h8 == readAddr[4:0] ? $signed(io_array_8) : $signed(_GEN_114); // @[AXIWrapperChiselInsertSort.scala 248:{22,22}]
  wire [7:0] _GEN_116 = 5'h9 == readAddr[4:0] ? $signed(io_array_9) : $signed(_GEN_115); // @[AXIWrapperChiselInsertSort.scala 248:{22,22}]
  wire [7:0] _GEN_117 = 5'ha == readAddr[4:0] ? $signed(io_array_10) : $signed(_GEN_116); // @[AXIWrapperChiselInsertSort.scala 248:{22,22}]
  wire [7:0] _GEN_118 = 5'hb == readAddr[4:0] ? $signed(io_array_11) : $signed(_GEN_117); // @[AXIWrapperChiselInsertSort.scala 248:{22,22}]
  wire [7:0] _GEN_119 = 5'hc == readAddr[4:0] ? $signed(io_array_12) : $signed(_GEN_118); // @[AXIWrapperChiselInsertSort.scala 248:{22,22}]
  wire [7:0] _GEN_120 = 5'hd == readAddr[4:0] ? $signed(io_array_13) : $signed(_GEN_119); // @[AXIWrapperChiselInsertSort.scala 248:{22,22}]
  wire [7:0] _GEN_121 = 5'he == readAddr[4:0] ? $signed(io_array_14) : $signed(_GEN_120); // @[AXIWrapperChiselInsertSort.scala 248:{22,22}]
  wire [7:0] _GEN_122 = 5'hf == readAddr[4:0] ? $signed(io_array_15) : $signed(_GEN_121); // @[AXIWrapperChiselInsertSort.scala 248:{22,22}]
  wire [7:0] _GEN_123 = 5'h10 == readAddr[4:0] ? $signed(io_array_16) : $signed(_GEN_122); // @[AXIWrapperChiselInsertSort.scala 248:{22,22}]
  wire [7:0] _GEN_124 = 5'h11 == readAddr[4:0] ? $signed(io_array_17) : $signed(_GEN_123); // @[AXIWrapperChiselInsertSort.scala 248:{22,22}]
  wire [7:0] _GEN_125 = 5'h12 == readAddr[4:0] ? $signed(io_array_18) : $signed(_GEN_124); // @[AXIWrapperChiselInsertSort.scala 248:{22,22}]
  wire [7:0] _GEN_126 = 5'h13 == readAddr[4:0] ? $signed(io_array_19) : $signed(_GEN_125); // @[AXIWrapperChiselInsertSort.scala 248:{22,22}]
  wire [7:0] _reg_data_out_T_2 = readAddr - 8'h14; // @[AXIWrapperChiselInsertSort.scala 250:47]
  wire [7:0] io_array_out_0 = modInsertSort_io_array_out_0[7:0]; // @[AXIWrapperChiselInsertSort.scala 232:25 71:28]
  wire [7:0] io_array_out_1 = modInsertSort_io_array_out_1[7:0]; // @[AXIWrapperChiselInsertSort.scala 232:25 71:28]
  wire [7:0] _GEN_128 = 5'h1 == _reg_data_out_T_2[4:0] ? $signed(io_array_out_1) : $signed(io_array_out_0); // @[AXIWrapperChiselInsertSort.scala 250:{22,22}]
  wire [7:0] io_array_out_2 = modInsertSort_io_array_out_2[7:0]; // @[AXIWrapperChiselInsertSort.scala 232:25 71:28]
  wire [7:0] _GEN_129 = 5'h2 == _reg_data_out_T_2[4:0] ? $signed(io_array_out_2) : $signed(_GEN_128); // @[AXIWrapperChiselInsertSort.scala 250:{22,22}]
  wire [7:0] io_array_out_3 = modInsertSort_io_array_out_3[7:0]; // @[AXIWrapperChiselInsertSort.scala 232:25 71:28]
  wire [7:0] _GEN_130 = 5'h3 == _reg_data_out_T_2[4:0] ? $signed(io_array_out_3) : $signed(_GEN_129); // @[AXIWrapperChiselInsertSort.scala 250:{22,22}]
  wire [7:0] io_array_out_4 = modInsertSort_io_array_out_4[7:0]; // @[AXIWrapperChiselInsertSort.scala 232:25 71:28]
  wire [7:0] _GEN_131 = 5'h4 == _reg_data_out_T_2[4:0] ? $signed(io_array_out_4) : $signed(_GEN_130); // @[AXIWrapperChiselInsertSort.scala 250:{22,22}]
  wire [7:0] io_array_out_5 = modInsertSort_io_array_out_5[7:0]; // @[AXIWrapperChiselInsertSort.scala 232:25 71:28]
  wire [7:0] _GEN_132 = 5'h5 == _reg_data_out_T_2[4:0] ? $signed(io_array_out_5) : $signed(_GEN_131); // @[AXIWrapperChiselInsertSort.scala 250:{22,22}]
  wire [7:0] io_array_out_6 = modInsertSort_io_array_out_6[7:0]; // @[AXIWrapperChiselInsertSort.scala 232:25 71:28]
  wire [7:0] _GEN_133 = 5'h6 == _reg_data_out_T_2[4:0] ? $signed(io_array_out_6) : $signed(_GEN_132); // @[AXIWrapperChiselInsertSort.scala 250:{22,22}]
  wire [7:0] io_array_out_7 = modInsertSort_io_array_out_7[7:0]; // @[AXIWrapperChiselInsertSort.scala 232:25 71:28]
  wire [7:0] _GEN_134 = 5'h7 == _reg_data_out_T_2[4:0] ? $signed(io_array_out_7) : $signed(_GEN_133); // @[AXIWrapperChiselInsertSort.scala 250:{22,22}]
  wire [7:0] io_array_out_8 = modInsertSort_io_array_out_8[7:0]; // @[AXIWrapperChiselInsertSort.scala 232:25 71:28]
  wire [7:0] _GEN_135 = 5'h8 == _reg_data_out_T_2[4:0] ? $signed(io_array_out_8) : $signed(_GEN_134); // @[AXIWrapperChiselInsertSort.scala 250:{22,22}]
  wire [7:0] io_array_out_9 = modInsertSort_io_array_out_9[7:0]; // @[AXIWrapperChiselInsertSort.scala 232:25 71:28]
  wire [7:0] _GEN_136 = 5'h9 == _reg_data_out_T_2[4:0] ? $signed(io_array_out_9) : $signed(_GEN_135); // @[AXIWrapperChiselInsertSort.scala 250:{22,22}]
  wire [7:0] io_array_out_10 = modInsertSort_io_array_out_10[7:0]; // @[AXIWrapperChiselInsertSort.scala 232:25 71:28]
  wire [7:0] _GEN_137 = 5'ha == _reg_data_out_T_2[4:0] ? $signed(io_array_out_10) : $signed(_GEN_136); // @[AXIWrapperChiselInsertSort.scala 250:{22,22}]
  wire [7:0] io_array_out_11 = modInsertSort_io_array_out_11[7:0]; // @[AXIWrapperChiselInsertSort.scala 232:25 71:28]
  wire [7:0] _GEN_138 = 5'hb == _reg_data_out_T_2[4:0] ? $signed(io_array_out_11) : $signed(_GEN_137); // @[AXIWrapperChiselInsertSort.scala 250:{22,22}]
  wire [7:0] io_array_out_12 = modInsertSort_io_array_out_12[7:0]; // @[AXIWrapperChiselInsertSort.scala 232:25 71:28]
  wire [7:0] _GEN_139 = 5'hc == _reg_data_out_T_2[4:0] ? $signed(io_array_out_12) : $signed(_GEN_138); // @[AXIWrapperChiselInsertSort.scala 250:{22,22}]
  wire [7:0] io_array_out_13 = modInsertSort_io_array_out_13[7:0]; // @[AXIWrapperChiselInsertSort.scala 232:25 71:28]
  wire [7:0] _GEN_140 = 5'hd == _reg_data_out_T_2[4:0] ? $signed(io_array_out_13) : $signed(_GEN_139); // @[AXIWrapperChiselInsertSort.scala 250:{22,22}]
  wire [7:0] io_array_out_14 = modInsertSort_io_array_out_14[7:0]; // @[AXIWrapperChiselInsertSort.scala 232:25 71:28]
  wire [7:0] _GEN_141 = 5'he == _reg_data_out_T_2[4:0] ? $signed(io_array_out_14) : $signed(_GEN_140); // @[AXIWrapperChiselInsertSort.scala 250:{22,22}]
  wire [7:0] io_array_out_15 = modInsertSort_io_array_out_15[7:0]; // @[AXIWrapperChiselInsertSort.scala 232:25 71:28]
  wire [7:0] _GEN_142 = 5'hf == _reg_data_out_T_2[4:0] ? $signed(io_array_out_15) : $signed(_GEN_141); // @[AXIWrapperChiselInsertSort.scala 250:{22,22}]
  wire [7:0] io_array_out_16 = modInsertSort_io_array_out_16[7:0]; // @[AXIWrapperChiselInsertSort.scala 232:25 71:28]
  wire [7:0] _GEN_143 = 5'h10 == _reg_data_out_T_2[4:0] ? $signed(io_array_out_16) : $signed(_GEN_142); // @[AXIWrapperChiselInsertSort.scala 250:{22,22}]
  wire [7:0] io_array_out_17 = modInsertSort_io_array_out_17[7:0]; // @[AXIWrapperChiselInsertSort.scala 232:25 71:28]
  wire [7:0] _GEN_144 = 5'h11 == _reg_data_out_T_2[4:0] ? $signed(io_array_out_17) : $signed(_GEN_143); // @[AXIWrapperChiselInsertSort.scala 250:{22,22}]
  wire [7:0] io_array_out_18 = modInsertSort_io_array_out_18[7:0]; // @[AXIWrapperChiselInsertSort.scala 232:25 71:28]
  wire [7:0] _GEN_145 = 5'h12 == _reg_data_out_T_2[4:0] ? $signed(io_array_out_18) : $signed(_GEN_144); // @[AXIWrapperChiselInsertSort.scala 250:{22,22}]
  wire [7:0] io_array_out_19 = modInsertSort_io_array_out_19[7:0]; // @[AXIWrapperChiselInsertSort.scala 232:25 71:28]
  wire [7:0] _GEN_146 = 5'h13 == _reg_data_out_T_2[4:0] ? $signed(io_array_out_19) : $signed(_GEN_145); // @[AXIWrapperChiselInsertSort.scala 250:{22,22}]
  wire [1:0] _reg_data_out_T_5 = {1'h0,io_ready}; // @[AXIWrapperChiselInsertSort.scala 254:44]
  wire [1:0] _GEN_147 = 8'h29 == readAddr ? $signed(_reg_data_out_T_5) : $signed(2'sh0); // @[AXIWrapperChiselInsertSort.scala 253:38 254:22 256:22]
  insertSort modInsertSort ( // @[AXIWrapperChiselInsertSort.scala 40:31]
    .clock(modInsertSort_clock),
    .reset(modInsertSort_reset),
    .io_array_0(modInsertSort_io_array_0),
    .io_array_1(modInsertSort_io_array_1),
    .io_array_2(modInsertSort_io_array_2),
    .io_array_3(modInsertSort_io_array_3),
    .io_array_4(modInsertSort_io_array_4),
    .io_array_5(modInsertSort_io_array_5),
    .io_array_6(modInsertSort_io_array_6),
    .io_array_7(modInsertSort_io_array_7),
    .io_array_8(modInsertSort_io_array_8),
    .io_array_9(modInsertSort_io_array_9),
    .io_array_10(modInsertSort_io_array_10),
    .io_array_11(modInsertSort_io_array_11),
    .io_array_12(modInsertSort_io_array_12),
    .io_array_13(modInsertSort_io_array_13),
    .io_array_14(modInsertSort_io_array_14),
    .io_array_15(modInsertSort_io_array_15),
    .io_array_16(modInsertSort_io_array_16),
    .io_array_17(modInsertSort_io_array_17),
    .io_array_18(modInsertSort_io_array_18),
    .io_array_19(modInsertSort_io_array_19),
    .io_valid(modInsertSort_io_valid),
    .io_array_out_0(modInsertSort_io_array_out_0),
    .io_array_out_1(modInsertSort_io_array_out_1),
    .io_array_out_2(modInsertSort_io_array_out_2),
    .io_array_out_3(modInsertSort_io_array_out_3),
    .io_array_out_4(modInsertSort_io_array_out_4),
    .io_array_out_5(modInsertSort_io_array_out_5),
    .io_array_out_6(modInsertSort_io_array_out_6),
    .io_array_out_7(modInsertSort_io_array_out_7),
    .io_array_out_8(modInsertSort_io_array_out_8),
    .io_array_out_9(modInsertSort_io_array_out_9),
    .io_array_out_10(modInsertSort_io_array_out_10),
    .io_array_out_11(modInsertSort_io_array_out_11),
    .io_array_out_12(modInsertSort_io_array_out_12),
    .io_array_out_13(modInsertSort_io_array_out_13),
    .io_array_out_14(modInsertSort_io_array_out_14),
    .io_array_out_15(modInsertSort_io_array_out_15),
    .io_array_out_16(modInsertSort_io_array_out_16),
    .io_array_out_17(modInsertSort_io_array_out_17),
    .io_array_out_18(modInsertSort_io_array_out_18),
    .io_array_out_19(modInsertSort_io_array_out_19),
    .io_ready(modInsertSort_io_ready)
  );
  assign io_S_AXI_AWREADY = axi_awready; // @[AXIWrapperChiselInsertSort.scala 78:22]
  assign io_S_AXI_WREADY = axi_wready; // @[AXIWrapperChiselInsertSort.scala 79:22]
  assign io_S_AXI_BRESP = 2'h0; // @[AXIWrapperChiselInsertSort.scala 80:22]
  assign io_S_AXI_BVALID = axi_bvalid; // @[AXIWrapperChiselInsertSort.scala 81:26]
  assign io_S_AXI_ARREADY = axi_arready; // @[AXIWrapperChiselInsertSort.scala 82:22]
  assign io_S_AXI_RDATA = axi_rdata; // @[AXIWrapperChiselInsertSort.scala 83:22]
  assign io_S_AXI_RRESP = 2'h0; // @[AXIWrapperChiselInsertSort.scala 84:22]
  assign io_S_AXI_RVALID = axi_rvalid; // @[AXIWrapperChiselInsertSort.scala 85:22]
  assign modInsertSort_clock = clock; // @[AXIWrapperChiselInsertSort.scala 221:25]
  assign modInsertSort_reset = reset; // @[AXIWrapperChiselInsertSort.scala 222:25]
  assign modInsertSort_io_array_0 = {{24{io_array_0[7]}},io_array_0}; // @[AXIWrapperChiselInsertSort.scala 227:39]
  assign modInsertSort_io_array_1 = {{24{io_array_1[7]}},io_array_1}; // @[AXIWrapperChiselInsertSort.scala 227:39]
  assign modInsertSort_io_array_2 = {{24{io_array_2[7]}},io_array_2}; // @[AXIWrapperChiselInsertSort.scala 227:39]
  assign modInsertSort_io_array_3 = {{24{io_array_3[7]}},io_array_3}; // @[AXIWrapperChiselInsertSort.scala 227:39]
  assign modInsertSort_io_array_4 = {{24{io_array_4[7]}},io_array_4}; // @[AXIWrapperChiselInsertSort.scala 227:39]
  assign modInsertSort_io_array_5 = {{24{io_array_5[7]}},io_array_5}; // @[AXIWrapperChiselInsertSort.scala 227:39]
  assign modInsertSort_io_array_6 = {{24{io_array_6[7]}},io_array_6}; // @[AXIWrapperChiselInsertSort.scala 227:39]
  assign modInsertSort_io_array_7 = {{24{io_array_7[7]}},io_array_7}; // @[AXIWrapperChiselInsertSort.scala 227:39]
  assign modInsertSort_io_array_8 = {{24{io_array_8[7]}},io_array_8}; // @[AXIWrapperChiselInsertSort.scala 227:39]
  assign modInsertSort_io_array_9 = {{24{io_array_9[7]}},io_array_9}; // @[AXIWrapperChiselInsertSort.scala 227:39]
  assign modInsertSort_io_array_10 = {{24{io_array_10[7]}},io_array_10}; // @[AXIWrapperChiselInsertSort.scala 227:39]
  assign modInsertSort_io_array_11 = {{24{io_array_11[7]}},io_array_11}; // @[AXIWrapperChiselInsertSort.scala 227:39]
  assign modInsertSort_io_array_12 = {{24{io_array_12[7]}},io_array_12}; // @[AXIWrapperChiselInsertSort.scala 227:39]
  assign modInsertSort_io_array_13 = {{24{io_array_13[7]}},io_array_13}; // @[AXIWrapperChiselInsertSort.scala 227:39]
  assign modInsertSort_io_array_14 = {{24{io_array_14[7]}},io_array_14}; // @[AXIWrapperChiselInsertSort.scala 227:39]
  assign modInsertSort_io_array_15 = {{24{io_array_15[7]}},io_array_15}; // @[AXIWrapperChiselInsertSort.scala 227:39]
  assign modInsertSort_io_array_16 = {{24{io_array_16[7]}},io_array_16}; // @[AXIWrapperChiselInsertSort.scala 227:39]
  assign modInsertSort_io_array_17 = {{24{io_array_17[7]}},io_array_17}; // @[AXIWrapperChiselInsertSort.scala 227:39]
  assign modInsertSort_io_array_18 = {{24{io_array_18[7]}},io_array_18}; // @[AXIWrapperChiselInsertSort.scala 227:39]
  assign modInsertSort_io_array_19 = {{24{io_array_19[7]}},io_array_19}; // @[AXIWrapperChiselInsertSort.scala 227:39]
  assign modInsertSort_io_valid = io_valid_reg[0]; // @[AXIWrapperChiselInsertSort.scala 223:43]
  always @(posedge clock) begin
    if (reset) begin // @[AXIWrapperChiselInsertSort.scala 115:24]
      axi_awaddr <= 32'h0; // @[AXIWrapperChiselInsertSort.scala 116:20]
    end else if (_T_4) begin // @[AXIWrapperChiselInsertSort.scala 118:76]
      axi_awaddr <= io_S_AXI_AWADDR; // @[AXIWrapperChiselInsertSort.scala 119:24]
    end
    if (reset) begin // @[AXIWrapperChiselInsertSort.scala 187:24]
      axi_araddr <= 32'h0; // @[AXIWrapperChiselInsertSort.scala 189:21]
    end else if (~axi_arready & io_S_AXI_ARVALID) begin // @[AXIWrapperChiselInsertSort.scala 191:48]
      axi_araddr <= io_S_AXI_ARADDR; // @[AXIWrapperChiselInsertSort.scala 194:25]
    end
    if (reset) begin // @[AXIWrapperChiselInsertSort.scala 91:24]
      axi_awready <= 1'h0; // @[AXIWrapperChiselInsertSort.scala 92:21]
    end else begin
      axi_awready <= _T_4;
    end
    if (reset) begin // @[AXIWrapperChiselInsertSort.scala 127:24]
      axi_wready <= 1'h0; // @[AXIWrapperChiselInsertSort.scala 128:20]
    end else begin
      axi_wready <= _T_15;
    end
    if (reset) begin // @[AXIWrapperChiselInsertSort.scala 167:24]
      axi_bvalid <= 1'h0; // @[AXIWrapperChiselInsertSort.scala 168:20]
    end else begin
      axi_bvalid <= _GEN_93;
    end
    if (reset) begin // @[AXIWrapperChiselInsertSort.scala 187:24]
      axi_arready <= 1'h0; // @[AXIWrapperChiselInsertSort.scala 188:21]
    end else begin
      axi_arready <= _T_30;
    end
    if (reset) begin // @[AXIWrapperChiselInsertSort.scala 260:24]
      axi_rdata <= 32'sh0; // @[AXIWrapperChiselInsertSort.scala 261:19]
    end else if (_T_34) begin // @[AXIWrapperChiselInsertSort.scala 266:28]
      axi_rdata <= reg_data_out; // @[AXIWrapperChiselInsertSort.scala 267:23]
    end
    if (reset) begin // @[AXIWrapperChiselInsertSort.scala 208:24]
      axi_rvalid <= 1'h0; // @[AXIWrapperChiselInsertSort.scala 209:20]
    end else begin
      axi_rvalid <= _GEN_102;
    end
    if (reset) begin // @[AXIWrapperChiselInsertSort.scala 150:24]
      io_valid_reg <= 32'sh0; // @[AXIWrapperChiselInsertSort.scala 151:22]
    end else if (axi_awaddr[9:2] == 8'h28) begin // @[AXIWrapperChiselInsertSort.scala 153:77]
      io_valid_reg <= io_S_AXI_WDATA; // @[AXIWrapperChiselInsertSort.scala 154:26]
    end
    if (!(reset)) begin // @[AXIWrapperChiselInsertSort.scala 150:24]
      if (!(axi_awaddr[9:2] == 8'h28)) begin // @[AXIWrapperChiselInsertSort.scala 153:77]
        if (slv_reg_wren) begin // @[AXIWrapperChiselInsertSort.scala 156:32]
          if (5'h0 == axi_awaddr[6:2]) begin // @[AXIWrapperChiselInsertSort.scala 157:78]
            io_array_0 <= _io_array_T_20; // @[AXIWrapperChiselInsertSort.scala 157:78]
          end
        end
      end
    end
    if (!(reset)) begin // @[AXIWrapperChiselInsertSort.scala 150:24]
      if (!(axi_awaddr[9:2] == 8'h28)) begin // @[AXIWrapperChiselInsertSort.scala 153:77]
        if (slv_reg_wren) begin // @[AXIWrapperChiselInsertSort.scala 156:32]
          if (5'h1 == axi_awaddr[6:2]) begin // @[AXIWrapperChiselInsertSort.scala 157:78]
            io_array_1 <= _io_array_T_20; // @[AXIWrapperChiselInsertSort.scala 157:78]
          end
        end
      end
    end
    if (!(reset)) begin // @[AXIWrapperChiselInsertSort.scala 150:24]
      if (!(axi_awaddr[9:2] == 8'h28)) begin // @[AXIWrapperChiselInsertSort.scala 153:77]
        if (slv_reg_wren) begin // @[AXIWrapperChiselInsertSort.scala 156:32]
          if (5'h2 == axi_awaddr[6:2]) begin // @[AXIWrapperChiselInsertSort.scala 157:78]
            io_array_2 <= _io_array_T_20; // @[AXIWrapperChiselInsertSort.scala 157:78]
          end
        end
      end
    end
    if (!(reset)) begin // @[AXIWrapperChiselInsertSort.scala 150:24]
      if (!(axi_awaddr[9:2] == 8'h28)) begin // @[AXIWrapperChiselInsertSort.scala 153:77]
        if (slv_reg_wren) begin // @[AXIWrapperChiselInsertSort.scala 156:32]
          if (5'h3 == axi_awaddr[6:2]) begin // @[AXIWrapperChiselInsertSort.scala 157:78]
            io_array_3 <= _io_array_T_20; // @[AXIWrapperChiselInsertSort.scala 157:78]
          end
        end
      end
    end
    if (!(reset)) begin // @[AXIWrapperChiselInsertSort.scala 150:24]
      if (!(axi_awaddr[9:2] == 8'h28)) begin // @[AXIWrapperChiselInsertSort.scala 153:77]
        if (slv_reg_wren) begin // @[AXIWrapperChiselInsertSort.scala 156:32]
          if (5'h4 == axi_awaddr[6:2]) begin // @[AXIWrapperChiselInsertSort.scala 157:78]
            io_array_4 <= _io_array_T_20; // @[AXIWrapperChiselInsertSort.scala 157:78]
          end
        end
      end
    end
    if (!(reset)) begin // @[AXIWrapperChiselInsertSort.scala 150:24]
      if (!(axi_awaddr[9:2] == 8'h28)) begin // @[AXIWrapperChiselInsertSort.scala 153:77]
        if (slv_reg_wren) begin // @[AXIWrapperChiselInsertSort.scala 156:32]
          if (5'h5 == axi_awaddr[6:2]) begin // @[AXIWrapperChiselInsertSort.scala 157:78]
            io_array_5 <= _io_array_T_20; // @[AXIWrapperChiselInsertSort.scala 157:78]
          end
        end
      end
    end
    if (!(reset)) begin // @[AXIWrapperChiselInsertSort.scala 150:24]
      if (!(axi_awaddr[9:2] == 8'h28)) begin // @[AXIWrapperChiselInsertSort.scala 153:77]
        if (slv_reg_wren) begin // @[AXIWrapperChiselInsertSort.scala 156:32]
          if (5'h6 == axi_awaddr[6:2]) begin // @[AXIWrapperChiselInsertSort.scala 157:78]
            io_array_6 <= _io_array_T_20; // @[AXIWrapperChiselInsertSort.scala 157:78]
          end
        end
      end
    end
    if (!(reset)) begin // @[AXIWrapperChiselInsertSort.scala 150:24]
      if (!(axi_awaddr[9:2] == 8'h28)) begin // @[AXIWrapperChiselInsertSort.scala 153:77]
        if (slv_reg_wren) begin // @[AXIWrapperChiselInsertSort.scala 156:32]
          if (5'h7 == axi_awaddr[6:2]) begin // @[AXIWrapperChiselInsertSort.scala 157:78]
            io_array_7 <= _io_array_T_20; // @[AXIWrapperChiselInsertSort.scala 157:78]
          end
        end
      end
    end
    if (!(reset)) begin // @[AXIWrapperChiselInsertSort.scala 150:24]
      if (!(axi_awaddr[9:2] == 8'h28)) begin // @[AXIWrapperChiselInsertSort.scala 153:77]
        if (slv_reg_wren) begin // @[AXIWrapperChiselInsertSort.scala 156:32]
          if (5'h8 == axi_awaddr[6:2]) begin // @[AXIWrapperChiselInsertSort.scala 157:78]
            io_array_8 <= _io_array_T_20; // @[AXIWrapperChiselInsertSort.scala 157:78]
          end
        end
      end
    end
    if (!(reset)) begin // @[AXIWrapperChiselInsertSort.scala 150:24]
      if (!(axi_awaddr[9:2] == 8'h28)) begin // @[AXIWrapperChiselInsertSort.scala 153:77]
        if (slv_reg_wren) begin // @[AXIWrapperChiselInsertSort.scala 156:32]
          if (5'h9 == axi_awaddr[6:2]) begin // @[AXIWrapperChiselInsertSort.scala 157:78]
            io_array_9 <= _io_array_T_20; // @[AXIWrapperChiselInsertSort.scala 157:78]
          end
        end
      end
    end
    if (!(reset)) begin // @[AXIWrapperChiselInsertSort.scala 150:24]
      if (!(axi_awaddr[9:2] == 8'h28)) begin // @[AXIWrapperChiselInsertSort.scala 153:77]
        if (slv_reg_wren) begin // @[AXIWrapperChiselInsertSort.scala 156:32]
          if (5'ha == axi_awaddr[6:2]) begin // @[AXIWrapperChiselInsertSort.scala 157:78]
            io_array_10 <= _io_array_T_20; // @[AXIWrapperChiselInsertSort.scala 157:78]
          end
        end
      end
    end
    if (!(reset)) begin // @[AXIWrapperChiselInsertSort.scala 150:24]
      if (!(axi_awaddr[9:2] == 8'h28)) begin // @[AXIWrapperChiselInsertSort.scala 153:77]
        if (slv_reg_wren) begin // @[AXIWrapperChiselInsertSort.scala 156:32]
          if (5'hb == axi_awaddr[6:2]) begin // @[AXIWrapperChiselInsertSort.scala 157:78]
            io_array_11 <= _io_array_T_20; // @[AXIWrapperChiselInsertSort.scala 157:78]
          end
        end
      end
    end
    if (!(reset)) begin // @[AXIWrapperChiselInsertSort.scala 150:24]
      if (!(axi_awaddr[9:2] == 8'h28)) begin // @[AXIWrapperChiselInsertSort.scala 153:77]
        if (slv_reg_wren) begin // @[AXIWrapperChiselInsertSort.scala 156:32]
          if (5'hc == axi_awaddr[6:2]) begin // @[AXIWrapperChiselInsertSort.scala 157:78]
            io_array_12 <= _io_array_T_20; // @[AXIWrapperChiselInsertSort.scala 157:78]
          end
        end
      end
    end
    if (!(reset)) begin // @[AXIWrapperChiselInsertSort.scala 150:24]
      if (!(axi_awaddr[9:2] == 8'h28)) begin // @[AXIWrapperChiselInsertSort.scala 153:77]
        if (slv_reg_wren) begin // @[AXIWrapperChiselInsertSort.scala 156:32]
          if (5'hd == axi_awaddr[6:2]) begin // @[AXIWrapperChiselInsertSort.scala 157:78]
            io_array_13 <= _io_array_T_20; // @[AXIWrapperChiselInsertSort.scala 157:78]
          end
        end
      end
    end
    if (!(reset)) begin // @[AXIWrapperChiselInsertSort.scala 150:24]
      if (!(axi_awaddr[9:2] == 8'h28)) begin // @[AXIWrapperChiselInsertSort.scala 153:77]
        if (slv_reg_wren) begin // @[AXIWrapperChiselInsertSort.scala 156:32]
          if (5'he == axi_awaddr[6:2]) begin // @[AXIWrapperChiselInsertSort.scala 157:78]
            io_array_14 <= _io_array_T_20; // @[AXIWrapperChiselInsertSort.scala 157:78]
          end
        end
      end
    end
    if (!(reset)) begin // @[AXIWrapperChiselInsertSort.scala 150:24]
      if (!(axi_awaddr[9:2] == 8'h28)) begin // @[AXIWrapperChiselInsertSort.scala 153:77]
        if (slv_reg_wren) begin // @[AXIWrapperChiselInsertSort.scala 156:32]
          if (5'hf == axi_awaddr[6:2]) begin // @[AXIWrapperChiselInsertSort.scala 157:78]
            io_array_15 <= _io_array_T_20; // @[AXIWrapperChiselInsertSort.scala 157:78]
          end
        end
      end
    end
    if (!(reset)) begin // @[AXIWrapperChiselInsertSort.scala 150:24]
      if (!(axi_awaddr[9:2] == 8'h28)) begin // @[AXIWrapperChiselInsertSort.scala 153:77]
        if (slv_reg_wren) begin // @[AXIWrapperChiselInsertSort.scala 156:32]
          if (5'h10 == axi_awaddr[6:2]) begin // @[AXIWrapperChiselInsertSort.scala 157:78]
            io_array_16 <= _io_array_T_20; // @[AXIWrapperChiselInsertSort.scala 157:78]
          end
        end
      end
    end
    if (!(reset)) begin // @[AXIWrapperChiselInsertSort.scala 150:24]
      if (!(axi_awaddr[9:2] == 8'h28)) begin // @[AXIWrapperChiselInsertSort.scala 153:77]
        if (slv_reg_wren) begin // @[AXIWrapperChiselInsertSort.scala 156:32]
          if (5'h11 == axi_awaddr[6:2]) begin // @[AXIWrapperChiselInsertSort.scala 157:78]
            io_array_17 <= _io_array_T_20; // @[AXIWrapperChiselInsertSort.scala 157:78]
          end
        end
      end
    end
    if (!(reset)) begin // @[AXIWrapperChiselInsertSort.scala 150:24]
      if (!(axi_awaddr[9:2] == 8'h28)) begin // @[AXIWrapperChiselInsertSort.scala 153:77]
        if (slv_reg_wren) begin // @[AXIWrapperChiselInsertSort.scala 156:32]
          if (5'h12 == axi_awaddr[6:2]) begin // @[AXIWrapperChiselInsertSort.scala 157:78]
            io_array_18 <= _io_array_T_20; // @[AXIWrapperChiselInsertSort.scala 157:78]
          end
        end
      end
    end
    if (!(reset)) begin // @[AXIWrapperChiselInsertSort.scala 150:24]
      if (!(axi_awaddr[9:2] == 8'h28)) begin // @[AXIWrapperChiselInsertSort.scala 153:77]
        if (slv_reg_wren) begin // @[AXIWrapperChiselInsertSort.scala 156:32]
          if (5'h13 == axi_awaddr[6:2]) begin // @[AXIWrapperChiselInsertSort.scala 157:78]
            io_array_19 <= _io_array_T_20; // @[AXIWrapperChiselInsertSort.scala 157:78]
          end
        end
      end
    end
    if (readAddr <= 8'h13) begin // @[AXIWrapperChiselInsertSort.scala 247:51]
      reg_data_out <= {{24{_GEN_126[7]}},_GEN_126}; // @[AXIWrapperChiselInsertSort.scala 248:22]
    end else if (8'h14 <= readAddr & readAddr <= 8'h27) begin // @[AXIWrapperChiselInsertSort.scala 249:59]
      reg_data_out <= {{24{_GEN_146[7]}},_GEN_146}; // @[AXIWrapperChiselInsertSort.scala 250:22]
    end else if (8'h28 == readAddr) begin // @[AXIWrapperChiselInsertSort.scala 251:38]
      reg_data_out <= io_valid_reg; // @[AXIWrapperChiselInsertSort.scala 252:22]
    end else begin
      reg_data_out <= {{30{_GEN_147[1]}},_GEN_147};
    end
    aw_en <= reset | _GEN_3; // @[AXIWrapperChiselInsertSort.scala 91:24 93:21]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  axi_awaddr = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  axi_araddr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  axi_awready = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  axi_wready = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  axi_bvalid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  axi_arready = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  axi_rdata = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  axi_rvalid = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  io_valid_reg = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  io_array_0 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  io_array_1 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  io_array_2 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  io_array_3 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  io_array_4 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  io_array_5 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  io_array_6 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  io_array_7 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  io_array_8 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  io_array_9 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  io_array_10 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  io_array_11 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  io_array_12 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  io_array_13 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  io_array_14 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  io_array_15 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  io_array_16 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  io_array_17 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  io_array_18 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  io_array_19 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  reg_data_out = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  aw_en = _RAND_30[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

[success] Total time: 3 s, completed Jan 28, 2025, 1:06:11 PM
