module insertSort(
  input         clock,
  input         reset,
  input  [31:0] io_array_0,
  input  [31:0] io_array_1,
  input  [31:0] io_array_2,
  input  [31:0] io_array_3,
  input  [31:0] io_array_4,
  input  [31:0] io_array_5,
  input  [31:0] io_array_6,
  input  [31:0] io_array_7,
  input  [31:0] io_array_8,
  input  [31:0] io_array_9,
  input  [31:0] io_array_10,
  input  [31:0] io_array_11,
  input  [31:0] io_array_12,
  input  [31:0] io_array_13,
  input  [31:0] io_array_14,
  input  [31:0] io_array_15,
  input  [31:0] io_array_16,
  input  [31:0] io_array_17,
  input  [31:0] io_array_18,
  input  [31:0] io_array_19,
  input         io_valid,
  output [31:0] io_array_out_0,
  output [31:0] io_array_out_1,
  output [31:0] io_array_out_2,
  output [31:0] io_array_out_3,
  output [31:0] io_array_out_4,
  output [31:0] io_array_out_5,
  output [31:0] io_array_out_6,
  output [31:0] io_array_out_7,
  output [31:0] io_array_out_8,
  output [31:0] io_array_out_9,
  output [31:0] io_array_out_10,
  output [31:0] io_array_out_11,
  output [31:0] io_array_out_12,
  output [31:0] io_array_out_13,
  output [31:0] io_array_out_14,
  output [31:0] io_array_out_15,
  output [31:0] io_array_out_16,
  output [31:0] io_array_out_17,
  output [31:0] io_array_out_18,
  output [31:0] io_array_out_19,
  output        io_ready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] state; // @[insertSort.scala 13:24]
  reg [31:0] array_0; // @[insertSort.scala 15:20]
  reg [31:0] array_1; // @[insertSort.scala 15:20]
  reg [31:0] array_2; // @[insertSort.scala 15:20]
  reg [31:0] array_3; // @[insertSort.scala 15:20]
  reg [31:0] array_4; // @[insertSort.scala 15:20]
  reg [31:0] array_5; // @[insertSort.scala 15:20]
  reg [31:0] array_6; // @[insertSort.scala 15:20]
  reg [31:0] array_7; // @[insertSort.scala 15:20]
  reg [31:0] array_8; // @[insertSort.scala 15:20]
  reg [31:0] array_9; // @[insertSort.scala 15:20]
  reg [31:0] array_10; // @[insertSort.scala 15:20]
  reg [31:0] array_11; // @[insertSort.scala 15:20]
  reg [31:0] array_12; // @[insertSort.scala 15:20]
  reg [31:0] array_13; // @[insertSort.scala 15:20]
  reg [31:0] array_14; // @[insertSort.scala 15:20]
  reg [31:0] array_15; // @[insertSort.scala 15:20]
  reg [31:0] array_16; // @[insertSort.scala 15:20]
  reg [31:0] array_17; // @[insertSort.scala 15:20]
  reg [31:0] array_18; // @[insertSort.scala 15:20]
  reg [31:0] array_19; // @[insertSort.scala 15:20]
  reg  REG; // @[insertSort.scala 16:17]
  wire [31:0] _GEN_0 = REG ? $signed(io_array_0) : $signed(array_0); // @[insertSort.scala 16:29 17:15 15:20]
  wire [31:0] _GEN_1 = REG ? $signed(io_array_1) : $signed(array_1); // @[insertSort.scala 16:29 17:15 15:20]
  wire [31:0] _GEN_2 = REG ? $signed(io_array_2) : $signed(array_2); // @[insertSort.scala 16:29 17:15 15:20]
  wire [31:0] _GEN_3 = REG ? $signed(io_array_3) : $signed(array_3); // @[insertSort.scala 16:29 17:15 15:20]
  wire [31:0] _GEN_4 = REG ? $signed(io_array_4) : $signed(array_4); // @[insertSort.scala 16:29 17:15 15:20]
  wire [31:0] _GEN_5 = REG ? $signed(io_array_5) : $signed(array_5); // @[insertSort.scala 16:29 17:15 15:20]
  wire [31:0] _GEN_6 = REG ? $signed(io_array_6) : $signed(array_6); // @[insertSort.scala 16:29 17:15 15:20]
  wire [31:0] _GEN_7 = REG ? $signed(io_array_7) : $signed(array_7); // @[insertSort.scala 16:29 17:15 15:20]
  wire [31:0] _GEN_8 = REG ? $signed(io_array_8) : $signed(array_8); // @[insertSort.scala 16:29 17:15 15:20]
  wire [31:0] _GEN_9 = REG ? $signed(io_array_9) : $signed(array_9); // @[insertSort.scala 16:29 17:15 15:20]
  wire [31:0] _GEN_10 = REG ? $signed(io_array_10) : $signed(array_10); // @[insertSort.scala 16:29 17:15 15:20]
  wire [31:0] _GEN_11 = REG ? $signed(io_array_11) : $signed(array_11); // @[insertSort.scala 16:29 17:15 15:20]
  wire [31:0] _GEN_12 = REG ? $signed(io_array_12) : $signed(array_12); // @[insertSort.scala 16:29 17:15 15:20]
  wire [31:0] _GEN_13 = REG ? $signed(io_array_13) : $signed(array_13); // @[insertSort.scala 16:29 17:15 15:20]
  wire [31:0] _GEN_14 = REG ? $signed(io_array_14) : $signed(array_14); // @[insertSort.scala 16:29 17:15 15:20]
  wire [31:0] _GEN_15 = REG ? $signed(io_array_15) : $signed(array_15); // @[insertSort.scala 16:29 17:15 15:20]
  wire [31:0] _GEN_16 = REG ? $signed(io_array_16) : $signed(array_16); // @[insertSort.scala 16:29 17:15 15:20]
  wire [31:0] _GEN_17 = REG ? $signed(io_array_17) : $signed(array_17); // @[insertSort.scala 16:29 17:15 15:20]
  wire [31:0] _GEN_18 = REG ? $signed(io_array_18) : $signed(array_18); // @[insertSort.scala 16:29 17:15 15:20]
  wire [31:0] _GEN_19 = REG ? $signed(io_array_19) : $signed(array_19); // @[insertSort.scala 16:29 17:15 15:20]
  reg [31:0] i; // @[insertSort.scala 20:16]
  reg [31:0] key; // @[insertSort.scala 21:18]
  reg [31:0] j; // @[insertSort.scala 22:16]
  wire [3:0] _state_T_2 = $signed(i) < 32'sha ? 4'h2 : 4'hc; // @[insertSort.scala 33:25]
  wire [31:0] _key_T = i; // @[insertSort.scala 36:36]
  wire [31:0] _GEN_21 = 5'h1 == _key_T[4:0] ? $signed(array_1) : $signed(array_0); // @[insertSort.scala 36:{17,17}]
  wire [31:0] _GEN_22 = 5'h2 == _key_T[4:0] ? $signed(array_2) : $signed(_GEN_21); // @[insertSort.scala 36:{17,17}]
  wire [31:0] _GEN_23 = 5'h3 == _key_T[4:0] ? $signed(array_3) : $signed(_GEN_22); // @[insertSort.scala 36:{17,17}]
  wire [31:0] _GEN_24 = 5'h4 == _key_T[4:0] ? $signed(array_4) : $signed(_GEN_23); // @[insertSort.scala 36:{17,17}]
  wire [31:0] _GEN_25 = 5'h5 == _key_T[4:0] ? $signed(array_5) : $signed(_GEN_24); // @[insertSort.scala 36:{17,17}]
  wire [31:0] _GEN_26 = 5'h6 == _key_T[4:0] ? $signed(array_6) : $signed(_GEN_25); // @[insertSort.scala 36:{17,17}]
  wire [31:0] _GEN_27 = 5'h7 == _key_T[4:0] ? $signed(array_7) : $signed(_GEN_26); // @[insertSort.scala 36:{17,17}]
  wire [31:0] _GEN_28 = 5'h8 == _key_T[4:0] ? $signed(array_8) : $signed(_GEN_27); // @[insertSort.scala 36:{17,17}]
  wire [31:0] _GEN_29 = 5'h9 == _key_T[4:0] ? $signed(array_9) : $signed(_GEN_28); // @[insertSort.scala 36:{17,17}]
  wire [31:0] _GEN_30 = 5'ha == _key_T[4:0] ? $signed(array_10) : $signed(_GEN_29); // @[insertSort.scala 36:{17,17}]
  wire [31:0] _GEN_31 = 5'hb == _key_T[4:0] ? $signed(array_11) : $signed(_GEN_30); // @[insertSort.scala 36:{17,17}]
  wire [31:0] _GEN_32 = 5'hc == _key_T[4:0] ? $signed(array_12) : $signed(_GEN_31); // @[insertSort.scala 36:{17,17}]
  wire [31:0] _GEN_33 = 5'hd == _key_T[4:0] ? $signed(array_13) : $signed(_GEN_32); // @[insertSort.scala 36:{17,17}]
  wire [31:0] _GEN_34 = 5'he == _key_T[4:0] ? $signed(array_14) : $signed(_GEN_33); // @[insertSort.scala 36:{17,17}]
  wire [31:0] _GEN_35 = 5'hf == _key_T[4:0] ? $signed(array_15) : $signed(_GEN_34); // @[insertSort.scala 36:{17,17}]
  wire [31:0] _GEN_36 = 5'h10 == _key_T[4:0] ? $signed(array_16) : $signed(_GEN_35); // @[insertSort.scala 36:{17,17}]
  wire [31:0] _GEN_37 = 5'h11 == _key_T[4:0] ? $signed(array_17) : $signed(_GEN_36); // @[insertSort.scala 36:{17,17}]
  wire [31:0] _GEN_38 = 5'h12 == _key_T[4:0] ? $signed(array_18) : $signed(_GEN_37); // @[insertSort.scala 36:{17,17}]
  wire [31:0] _GEN_39 = 5'h13 == _key_T[4:0] ? $signed(array_19) : $signed(_GEN_38); // @[insertSort.scala 36:{17,17}]
  wire [31:0] _j_T_2 = $signed(i) - 32'sh1; // @[insertSort.scala 40:20]
  wire [31:0] _state_T_4 = j; // @[insertSort.scala 44:54]
  wire [31:0] _GEN_41 = 5'h1 == _state_T_4[4:0] ? $signed(array_1) : $signed(array_0); // @[insertSort.scala 44:{58,58}]
  wire [31:0] _GEN_42 = 5'h2 == _state_T_4[4:0] ? $signed(array_2) : $signed(_GEN_41); // @[insertSort.scala 44:{58,58}]
  wire [31:0] _GEN_43 = 5'h3 == _state_T_4[4:0] ? $signed(array_3) : $signed(_GEN_42); // @[insertSort.scala 44:{58,58}]
  wire [31:0] _GEN_44 = 5'h4 == _state_T_4[4:0] ? $signed(array_4) : $signed(_GEN_43); // @[insertSort.scala 44:{58,58}]
  wire [31:0] _GEN_45 = 5'h5 == _state_T_4[4:0] ? $signed(array_5) : $signed(_GEN_44); // @[insertSort.scala 44:{58,58}]
  wire [31:0] _GEN_46 = 5'h6 == _state_T_4[4:0] ? $signed(array_6) : $signed(_GEN_45); // @[insertSort.scala 44:{58,58}]
  wire [31:0] _GEN_47 = 5'h7 == _state_T_4[4:0] ? $signed(array_7) : $signed(_GEN_46); // @[insertSort.scala 44:{58,58}]
  wire [31:0] _GEN_48 = 5'h8 == _state_T_4[4:0] ? $signed(array_8) : $signed(_GEN_47); // @[insertSort.scala 44:{58,58}]
  wire [31:0] _GEN_49 = 5'h9 == _state_T_4[4:0] ? $signed(array_9) : $signed(_GEN_48); // @[insertSort.scala 44:{58,58}]
  wire [31:0] _GEN_50 = 5'ha == _state_T_4[4:0] ? $signed(array_10) : $signed(_GEN_49); // @[insertSort.scala 44:{58,58}]
  wire [31:0] _GEN_51 = 5'hb == _state_T_4[4:0] ? $signed(array_11) : $signed(_GEN_50); // @[insertSort.scala 44:{58,58}]
  wire [31:0] _GEN_52 = 5'hc == _state_T_4[4:0] ? $signed(array_12) : $signed(_GEN_51); // @[insertSort.scala 44:{58,58}]
  wire [31:0] _GEN_53 = 5'hd == _state_T_4[4:0] ? $signed(array_13) : $signed(_GEN_52); // @[insertSort.scala 44:{58,58}]
  wire [31:0] _GEN_54 = 5'he == _state_T_4[4:0] ? $signed(array_14) : $signed(_GEN_53); // @[insertSort.scala 44:{58,58}]
  wire [31:0] _GEN_55 = 5'hf == _state_T_4[4:0] ? $signed(array_15) : $signed(_GEN_54); // @[insertSort.scala 44:{58,58}]
  wire [31:0] _GEN_56 = 5'h10 == _state_T_4[4:0] ? $signed(array_16) : $signed(_GEN_55); // @[insertSort.scala 44:{58,58}]
  wire [31:0] _GEN_57 = 5'h11 == _state_T_4[4:0] ? $signed(array_17) : $signed(_GEN_56); // @[insertSort.scala 44:{58,58}]
  wire [31:0] _GEN_58 = 5'h12 == _state_T_4[4:0] ? $signed(array_18) : $signed(_GEN_57); // @[insertSort.scala 44:{58,58}]
  wire [31:0] _GEN_59 = 5'h13 == _state_T_4[4:0] ? $signed(array_19) : $signed(_GEN_58); // @[insertSort.scala 44:{58,58}]
  wire  _state_T_6 = $signed(_GEN_59) > $signed(key); // @[insertSort.scala 44:58]
  wire [2:0] _state_T_8 = $signed(j) > 32'sh0 & $signed(_GEN_59) > $signed(key) ? 3'h5 : 3'h7; // @[insertSort.scala 44:25]
  wire [31:0] _T_11 = $signed(j) + 32'sh1; // @[insertSort.scala 47:36]
  wire [31:0] _GEN_60 = 5'h0 == _T_11[4:0] ? $signed(_GEN_59) : $signed(_GEN_0); // @[insertSort.scala 47:{40,40}]
  wire [31:0] _GEN_61 = 5'h1 == _T_11[4:0] ? $signed(_GEN_59) : $signed(_GEN_1); // @[insertSort.scala 47:{40,40}]
  wire [31:0] _GEN_62 = 5'h2 == _T_11[4:0] ? $signed(_GEN_59) : $signed(_GEN_2); // @[insertSort.scala 47:{40,40}]
  wire [31:0] _GEN_63 = 5'h3 == _T_11[4:0] ? $signed(_GEN_59) : $signed(_GEN_3); // @[insertSort.scala 47:{40,40}]
  wire [31:0] _GEN_64 = 5'h4 == _T_11[4:0] ? $signed(_GEN_59) : $signed(_GEN_4); // @[insertSort.scala 47:{40,40}]
  wire [31:0] _GEN_65 = 5'h5 == _T_11[4:0] ? $signed(_GEN_59) : $signed(_GEN_5); // @[insertSort.scala 47:{40,40}]
  wire [31:0] _GEN_66 = 5'h6 == _T_11[4:0] ? $signed(_GEN_59) : $signed(_GEN_6); // @[insertSort.scala 47:{40,40}]
  wire [31:0] _GEN_67 = 5'h7 == _T_11[4:0] ? $signed(_GEN_59) : $signed(_GEN_7); // @[insertSort.scala 47:{40,40}]
  wire [31:0] _GEN_68 = 5'h8 == _T_11[4:0] ? $signed(_GEN_59) : $signed(_GEN_8); // @[insertSort.scala 47:{40,40}]
  wire [31:0] _GEN_69 = 5'h9 == _T_11[4:0] ? $signed(_GEN_59) : $signed(_GEN_9); // @[insertSort.scala 47:{40,40}]
  wire [31:0] _GEN_70 = 5'ha == _T_11[4:0] ? $signed(_GEN_59) : $signed(_GEN_10); // @[insertSort.scala 47:{40,40}]
  wire [31:0] _GEN_71 = 5'hb == _T_11[4:0] ? $signed(_GEN_59) : $signed(_GEN_11); // @[insertSort.scala 47:{40,40}]
  wire [31:0] _GEN_72 = 5'hc == _T_11[4:0] ? $signed(_GEN_59) : $signed(_GEN_12); // @[insertSort.scala 47:{40,40}]
  wire [31:0] _GEN_73 = 5'hd == _T_11[4:0] ? $signed(_GEN_59) : $signed(_GEN_13); // @[insertSort.scala 47:{40,40}]
  wire [31:0] _GEN_74 = 5'he == _T_11[4:0] ? $signed(_GEN_59) : $signed(_GEN_14); // @[insertSort.scala 47:{40,40}]
  wire [31:0] _GEN_75 = 5'hf == _T_11[4:0] ? $signed(_GEN_59) : $signed(_GEN_15); // @[insertSort.scala 47:{40,40}]
  wire [31:0] _GEN_76 = 5'h10 == _T_11[4:0] ? $signed(_GEN_59) : $signed(_GEN_16); // @[insertSort.scala 47:{40,40}]
  wire [31:0] _GEN_77 = 5'h11 == _T_11[4:0] ? $signed(_GEN_59) : $signed(_GEN_17); // @[insertSort.scala 47:{40,40}]
  wire [31:0] _GEN_78 = 5'h12 == _T_11[4:0] ? $signed(_GEN_59) : $signed(_GEN_18); // @[insertSort.scala 47:{40,40}]
  wire [31:0] _GEN_79 = 5'h13 == _T_11[4:0] ? $signed(_GEN_59) : $signed(_GEN_19); // @[insertSort.scala 47:{40,40}]
  wire [31:0] _j_T_5 = $signed(j) - 32'sh1; // @[insertSort.scala 51:20]
  wire [3:0] _state_T_14 = $signed(j) == 32'sh0 & _state_T_6 ? 4'h8 : 4'ha; // @[insertSort.scala 55:25]
  wire [31:0] _GEN_160 = 5'h0 == _state_T_4[4:0] ? $signed(key) : $signed(_GEN_0); // @[insertSort.scala 62:{33,33}]
  wire [31:0] _GEN_161 = 5'h1 == _state_T_4[4:0] ? $signed(key) : $signed(_GEN_1); // @[insertSort.scala 62:{33,33}]
  wire [31:0] _GEN_162 = 5'h2 == _state_T_4[4:0] ? $signed(key) : $signed(_GEN_2); // @[insertSort.scala 62:{33,33}]
  wire [31:0] _GEN_163 = 5'h3 == _state_T_4[4:0] ? $signed(key) : $signed(_GEN_3); // @[insertSort.scala 62:{33,33}]
  wire [31:0] _GEN_164 = 5'h4 == _state_T_4[4:0] ? $signed(key) : $signed(_GEN_4); // @[insertSort.scala 62:{33,33}]
  wire [31:0] _GEN_165 = 5'h5 == _state_T_4[4:0] ? $signed(key) : $signed(_GEN_5); // @[insertSort.scala 62:{33,33}]
  wire [31:0] _GEN_166 = 5'h6 == _state_T_4[4:0] ? $signed(key) : $signed(_GEN_6); // @[insertSort.scala 62:{33,33}]
  wire [31:0] _GEN_167 = 5'h7 == _state_T_4[4:0] ? $signed(key) : $signed(_GEN_7); // @[insertSort.scala 62:{33,33}]
  wire [31:0] _GEN_168 = 5'h8 == _state_T_4[4:0] ? $signed(key) : $signed(_GEN_8); // @[insertSort.scala 62:{33,33}]
  wire [31:0] _GEN_169 = 5'h9 == _state_T_4[4:0] ? $signed(key) : $signed(_GEN_9); // @[insertSort.scala 62:{33,33}]
  wire [31:0] _GEN_170 = 5'ha == _state_T_4[4:0] ? $signed(key) : $signed(_GEN_10); // @[insertSort.scala 62:{33,33}]
  wire [31:0] _GEN_171 = 5'hb == _state_T_4[4:0] ? $signed(key) : $signed(_GEN_11); // @[insertSort.scala 62:{33,33}]
  wire [31:0] _GEN_172 = 5'hc == _state_T_4[4:0] ? $signed(key) : $signed(_GEN_12); // @[insertSort.scala 62:{33,33}]
  wire [31:0] _GEN_173 = 5'hd == _state_T_4[4:0] ? $signed(key) : $signed(_GEN_13); // @[insertSort.scala 62:{33,33}]
  wire [31:0] _GEN_174 = 5'he == _state_T_4[4:0] ? $signed(key) : $signed(_GEN_14); // @[insertSort.scala 62:{33,33}]
  wire [31:0] _GEN_175 = 5'hf == _state_T_4[4:0] ? $signed(key) : $signed(_GEN_15); // @[insertSort.scala 62:{33,33}]
  wire [31:0] _GEN_176 = 5'h10 == _state_T_4[4:0] ? $signed(key) : $signed(_GEN_16); // @[insertSort.scala 62:{33,33}]
  wire [31:0] _GEN_177 = 5'h11 == _state_T_4[4:0] ? $signed(key) : $signed(_GEN_17); // @[insertSort.scala 62:{33,33}]
  wire [31:0] _GEN_178 = 5'h12 == _state_T_4[4:0] ? $signed(key) : $signed(_GEN_18); // @[insertSort.scala 62:{33,33}]
  wire [31:0] _GEN_179 = 5'h13 == _state_T_4[4:0] ? $signed(key) : $signed(_GEN_19); // @[insertSort.scala 62:{33,33}]
  wire [31:0] _GEN_180 = 5'h0 == _T_11[4:0] ? $signed(key) : $signed(_GEN_0); // @[insertSort.scala 66:{40,40}]
  wire [31:0] _GEN_181 = 5'h1 == _T_11[4:0] ? $signed(key) : $signed(_GEN_1); // @[insertSort.scala 66:{40,40}]
  wire [31:0] _GEN_182 = 5'h2 == _T_11[4:0] ? $signed(key) : $signed(_GEN_2); // @[insertSort.scala 66:{40,40}]
  wire [31:0] _GEN_183 = 5'h3 == _T_11[4:0] ? $signed(key) : $signed(_GEN_3); // @[insertSort.scala 66:{40,40}]
  wire [31:0] _GEN_184 = 5'h4 == _T_11[4:0] ? $signed(key) : $signed(_GEN_4); // @[insertSort.scala 66:{40,40}]
  wire [31:0] _GEN_185 = 5'h5 == _T_11[4:0] ? $signed(key) : $signed(_GEN_5); // @[insertSort.scala 66:{40,40}]
  wire [31:0] _GEN_186 = 5'h6 == _T_11[4:0] ? $signed(key) : $signed(_GEN_6); // @[insertSort.scala 66:{40,40}]
  wire [31:0] _GEN_187 = 5'h7 == _T_11[4:0] ? $signed(key) : $signed(_GEN_7); // @[insertSort.scala 66:{40,40}]
  wire [31:0] _GEN_188 = 5'h8 == _T_11[4:0] ? $signed(key) : $signed(_GEN_8); // @[insertSort.scala 66:{40,40}]
  wire [31:0] _GEN_189 = 5'h9 == _T_11[4:0] ? $signed(key) : $signed(_GEN_9); // @[insertSort.scala 66:{40,40}]
  wire [31:0] _GEN_190 = 5'ha == _T_11[4:0] ? $signed(key) : $signed(_GEN_10); // @[insertSort.scala 66:{40,40}]
  wire [31:0] _GEN_191 = 5'hb == _T_11[4:0] ? $signed(key) : $signed(_GEN_11); // @[insertSort.scala 66:{40,40}]
  wire [31:0] _GEN_192 = 5'hc == _T_11[4:0] ? $signed(key) : $signed(_GEN_12); // @[insertSort.scala 66:{40,40}]
  wire [31:0] _GEN_193 = 5'hd == _T_11[4:0] ? $signed(key) : $signed(_GEN_13); // @[insertSort.scala 66:{40,40}]
  wire [31:0] _GEN_194 = 5'he == _T_11[4:0] ? $signed(key) : $signed(_GEN_14); // @[insertSort.scala 66:{40,40}]
  wire [31:0] _GEN_195 = 5'hf == _T_11[4:0] ? $signed(key) : $signed(_GEN_15); // @[insertSort.scala 66:{40,40}]
  wire [31:0] _GEN_196 = 5'h10 == _T_11[4:0] ? $signed(key) : $signed(_GEN_16); // @[insertSort.scala 66:{40,40}]
  wire [31:0] _GEN_197 = 5'h11 == _T_11[4:0] ? $signed(key) : $signed(_GEN_17); // @[insertSort.scala 66:{40,40}]
  wire [31:0] _GEN_198 = 5'h12 == _T_11[4:0] ? $signed(key) : $signed(_GEN_18); // @[insertSort.scala 66:{40,40}]
  wire [31:0] _GEN_199 = 5'h13 == _T_11[4:0] ? $signed(key) : $signed(_GEN_19); // @[insertSort.scala 66:{40,40}]
  wire [31:0] _i_T_2 = $signed(i) + 32'sh1; // @[insertSort.scala 70:21]
  wire [3:0] _GEN_200 = 4'hc == state ? 4'hf : state; // @[insertSort.scala 24:19 74:19 13:24]
  wire [31:0] _GEN_201 = 4'hb == state ? $signed(_i_T_2) : $signed(i); // @[insertSort.scala 24:19 70:15 20:16]
  wire [3:0] _GEN_202 = 4'hb == state ? 4'h1 : _GEN_200; // @[insertSort.scala 24:19 71:19]
  wire [31:0] _GEN_203 = 4'ha == state ? $signed(_GEN_180) : $signed(_GEN_0); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_204 = 4'ha == state ? $signed(_GEN_181) : $signed(_GEN_1); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_205 = 4'ha == state ? $signed(_GEN_182) : $signed(_GEN_2); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_206 = 4'ha == state ? $signed(_GEN_183) : $signed(_GEN_3); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_207 = 4'ha == state ? $signed(_GEN_184) : $signed(_GEN_4); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_208 = 4'ha == state ? $signed(_GEN_185) : $signed(_GEN_5); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_209 = 4'ha == state ? $signed(_GEN_186) : $signed(_GEN_6); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_210 = 4'ha == state ? $signed(_GEN_187) : $signed(_GEN_7); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_211 = 4'ha == state ? $signed(_GEN_188) : $signed(_GEN_8); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_212 = 4'ha == state ? $signed(_GEN_189) : $signed(_GEN_9); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_213 = 4'ha == state ? $signed(_GEN_190) : $signed(_GEN_10); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_214 = 4'ha == state ? $signed(_GEN_191) : $signed(_GEN_11); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_215 = 4'ha == state ? $signed(_GEN_192) : $signed(_GEN_12); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_216 = 4'ha == state ? $signed(_GEN_193) : $signed(_GEN_13); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_217 = 4'ha == state ? $signed(_GEN_194) : $signed(_GEN_14); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_218 = 4'ha == state ? $signed(_GEN_195) : $signed(_GEN_15); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_219 = 4'ha == state ? $signed(_GEN_196) : $signed(_GEN_16); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_220 = 4'ha == state ? $signed(_GEN_197) : $signed(_GEN_17); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_221 = 4'ha == state ? $signed(_GEN_198) : $signed(_GEN_18); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_222 = 4'ha == state ? $signed(_GEN_199) : $signed(_GEN_19); // @[insertSort.scala 24:19]
  wire [3:0] _GEN_223 = 4'ha == state ? 4'hb : _GEN_202; // @[insertSort.scala 24:19 67:19]
  wire [31:0] _GEN_224 = 4'ha == state ? $signed(i) : $signed(_GEN_201); // @[insertSort.scala 20:16 24:19]
  wire [31:0] _GEN_225 = 4'h9 == state ? $signed(_GEN_160) : $signed(_GEN_203); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_226 = 4'h9 == state ? $signed(_GEN_161) : $signed(_GEN_204); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_227 = 4'h9 == state ? $signed(_GEN_162) : $signed(_GEN_205); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_228 = 4'h9 == state ? $signed(_GEN_163) : $signed(_GEN_206); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_229 = 4'h9 == state ? $signed(_GEN_164) : $signed(_GEN_207); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_230 = 4'h9 == state ? $signed(_GEN_165) : $signed(_GEN_208); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_231 = 4'h9 == state ? $signed(_GEN_166) : $signed(_GEN_209); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_232 = 4'h9 == state ? $signed(_GEN_167) : $signed(_GEN_210); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_233 = 4'h9 == state ? $signed(_GEN_168) : $signed(_GEN_211); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_234 = 4'h9 == state ? $signed(_GEN_169) : $signed(_GEN_212); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_235 = 4'h9 == state ? $signed(_GEN_170) : $signed(_GEN_213); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_236 = 4'h9 == state ? $signed(_GEN_171) : $signed(_GEN_214); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_237 = 4'h9 == state ? $signed(_GEN_172) : $signed(_GEN_215); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_238 = 4'h9 == state ? $signed(_GEN_173) : $signed(_GEN_216); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_239 = 4'h9 == state ? $signed(_GEN_174) : $signed(_GEN_217); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_240 = 4'h9 == state ? $signed(_GEN_175) : $signed(_GEN_218); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_241 = 4'h9 == state ? $signed(_GEN_176) : $signed(_GEN_219); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_242 = 4'h9 == state ? $signed(_GEN_177) : $signed(_GEN_220); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_243 = 4'h9 == state ? $signed(_GEN_178) : $signed(_GEN_221); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_244 = 4'h9 == state ? $signed(_GEN_179) : $signed(_GEN_222); // @[insertSort.scala 24:19]
  wire [3:0] _GEN_245 = 4'h9 == state ? 4'hb : _GEN_223; // @[insertSort.scala 24:19 63:19]
  wire [31:0] _GEN_246 = 4'h9 == state ? $signed(i) : $signed(_GEN_224); // @[insertSort.scala 20:16 24:19]
  wire [31:0] _GEN_247 = 4'h8 == state ? $signed(_GEN_60) : $signed(_GEN_225); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_248 = 4'h8 == state ? $signed(_GEN_61) : $signed(_GEN_226); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_249 = 4'h8 == state ? $signed(_GEN_62) : $signed(_GEN_227); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_250 = 4'h8 == state ? $signed(_GEN_63) : $signed(_GEN_228); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_251 = 4'h8 == state ? $signed(_GEN_64) : $signed(_GEN_229); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_252 = 4'h8 == state ? $signed(_GEN_65) : $signed(_GEN_230); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_253 = 4'h8 == state ? $signed(_GEN_66) : $signed(_GEN_231); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_254 = 4'h8 == state ? $signed(_GEN_67) : $signed(_GEN_232); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_255 = 4'h8 == state ? $signed(_GEN_68) : $signed(_GEN_233); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_256 = 4'h8 == state ? $signed(_GEN_69) : $signed(_GEN_234); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_257 = 4'h8 == state ? $signed(_GEN_70) : $signed(_GEN_235); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_258 = 4'h8 == state ? $signed(_GEN_71) : $signed(_GEN_236); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_259 = 4'h8 == state ? $signed(_GEN_72) : $signed(_GEN_237); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_260 = 4'h8 == state ? $signed(_GEN_73) : $signed(_GEN_238); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_261 = 4'h8 == state ? $signed(_GEN_74) : $signed(_GEN_239); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_262 = 4'h8 == state ? $signed(_GEN_75) : $signed(_GEN_240); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_263 = 4'h8 == state ? $signed(_GEN_76) : $signed(_GEN_241); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_264 = 4'h8 == state ? $signed(_GEN_77) : $signed(_GEN_242); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_265 = 4'h8 == state ? $signed(_GEN_78) : $signed(_GEN_243); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_266 = 4'h8 == state ? $signed(_GEN_79) : $signed(_GEN_244); // @[insertSort.scala 24:19]
  wire [3:0] _GEN_267 = 4'h8 == state ? 4'h9 : _GEN_245; // @[insertSort.scala 24:19 59:19]
  wire [31:0] _GEN_268 = 4'h8 == state ? $signed(i) : $signed(_GEN_246); // @[insertSort.scala 20:16 24:19]
  wire [3:0] _GEN_269 = 4'h7 == state ? _state_T_14 : _GEN_267; // @[insertSort.scala 24:19 55:19]
  wire [31:0] _GEN_270 = 4'h7 == state ? $signed(_GEN_0) : $signed(_GEN_247); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_271 = 4'h7 == state ? $signed(_GEN_1) : $signed(_GEN_248); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_272 = 4'h7 == state ? $signed(_GEN_2) : $signed(_GEN_249); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_273 = 4'h7 == state ? $signed(_GEN_3) : $signed(_GEN_250); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_274 = 4'h7 == state ? $signed(_GEN_4) : $signed(_GEN_251); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_275 = 4'h7 == state ? $signed(_GEN_5) : $signed(_GEN_252); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_276 = 4'h7 == state ? $signed(_GEN_6) : $signed(_GEN_253); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_277 = 4'h7 == state ? $signed(_GEN_7) : $signed(_GEN_254); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_278 = 4'h7 == state ? $signed(_GEN_8) : $signed(_GEN_255); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_279 = 4'h7 == state ? $signed(_GEN_9) : $signed(_GEN_256); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_280 = 4'h7 == state ? $signed(_GEN_10) : $signed(_GEN_257); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_281 = 4'h7 == state ? $signed(_GEN_11) : $signed(_GEN_258); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_282 = 4'h7 == state ? $signed(_GEN_12) : $signed(_GEN_259); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_283 = 4'h7 == state ? $signed(_GEN_13) : $signed(_GEN_260); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_284 = 4'h7 == state ? $signed(_GEN_14) : $signed(_GEN_261); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_285 = 4'h7 == state ? $signed(_GEN_15) : $signed(_GEN_262); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_286 = 4'h7 == state ? $signed(_GEN_16) : $signed(_GEN_263); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_287 = 4'h7 == state ? $signed(_GEN_17) : $signed(_GEN_264); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_288 = 4'h7 == state ? $signed(_GEN_18) : $signed(_GEN_265); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_289 = 4'h7 == state ? $signed(_GEN_19) : $signed(_GEN_266); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_290 = 4'h7 == state ? $signed(i) : $signed(_GEN_268); // @[insertSort.scala 20:16 24:19]
  wire [31:0] _GEN_291 = 4'h6 == state ? $signed(_j_T_5) : $signed(j); // @[insertSort.scala 24:19 51:15 22:16]
  wire [3:0] _GEN_292 = 4'h6 == state ? 4'h4 : _GEN_269; // @[insertSort.scala 24:19 52:19]
  wire [31:0] _GEN_293 = 4'h6 == state ? $signed(_GEN_0) : $signed(_GEN_270); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_294 = 4'h6 == state ? $signed(_GEN_1) : $signed(_GEN_271); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_295 = 4'h6 == state ? $signed(_GEN_2) : $signed(_GEN_272); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_296 = 4'h6 == state ? $signed(_GEN_3) : $signed(_GEN_273); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_297 = 4'h6 == state ? $signed(_GEN_4) : $signed(_GEN_274); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_298 = 4'h6 == state ? $signed(_GEN_5) : $signed(_GEN_275); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_299 = 4'h6 == state ? $signed(_GEN_6) : $signed(_GEN_276); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_300 = 4'h6 == state ? $signed(_GEN_7) : $signed(_GEN_277); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_301 = 4'h6 == state ? $signed(_GEN_8) : $signed(_GEN_278); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_302 = 4'h6 == state ? $signed(_GEN_9) : $signed(_GEN_279); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_303 = 4'h6 == state ? $signed(_GEN_10) : $signed(_GEN_280); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_304 = 4'h6 == state ? $signed(_GEN_11) : $signed(_GEN_281); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_305 = 4'h6 == state ? $signed(_GEN_12) : $signed(_GEN_282); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_306 = 4'h6 == state ? $signed(_GEN_13) : $signed(_GEN_283); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_307 = 4'h6 == state ? $signed(_GEN_14) : $signed(_GEN_284); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_308 = 4'h6 == state ? $signed(_GEN_15) : $signed(_GEN_285); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_309 = 4'h6 == state ? $signed(_GEN_16) : $signed(_GEN_286); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_310 = 4'h6 == state ? $signed(_GEN_17) : $signed(_GEN_287); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_311 = 4'h6 == state ? $signed(_GEN_18) : $signed(_GEN_288); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_312 = 4'h6 == state ? $signed(_GEN_19) : $signed(_GEN_289); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_313 = 4'h6 == state ? $signed(i) : $signed(_GEN_290); // @[insertSort.scala 20:16 24:19]
  wire [31:0] _GEN_314 = 4'h5 == state ? $signed(_GEN_60) : $signed(_GEN_293); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_315 = 4'h5 == state ? $signed(_GEN_61) : $signed(_GEN_294); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_316 = 4'h5 == state ? $signed(_GEN_62) : $signed(_GEN_295); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_317 = 4'h5 == state ? $signed(_GEN_63) : $signed(_GEN_296); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_318 = 4'h5 == state ? $signed(_GEN_64) : $signed(_GEN_297); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_319 = 4'h5 == state ? $signed(_GEN_65) : $signed(_GEN_298); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_320 = 4'h5 == state ? $signed(_GEN_66) : $signed(_GEN_299); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_321 = 4'h5 == state ? $signed(_GEN_67) : $signed(_GEN_300); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_322 = 4'h5 == state ? $signed(_GEN_68) : $signed(_GEN_301); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_323 = 4'h5 == state ? $signed(_GEN_69) : $signed(_GEN_302); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_324 = 4'h5 == state ? $signed(_GEN_70) : $signed(_GEN_303); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_325 = 4'h5 == state ? $signed(_GEN_71) : $signed(_GEN_304); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_326 = 4'h5 == state ? $signed(_GEN_72) : $signed(_GEN_305); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_327 = 4'h5 == state ? $signed(_GEN_73) : $signed(_GEN_306); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_328 = 4'h5 == state ? $signed(_GEN_74) : $signed(_GEN_307); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_329 = 4'h5 == state ? $signed(_GEN_75) : $signed(_GEN_308); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_330 = 4'h5 == state ? $signed(_GEN_76) : $signed(_GEN_309); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_331 = 4'h5 == state ? $signed(_GEN_77) : $signed(_GEN_310); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_332 = 4'h5 == state ? $signed(_GEN_78) : $signed(_GEN_311); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_333 = 4'h5 == state ? $signed(_GEN_79) : $signed(_GEN_312); // @[insertSort.scala 24:19]
  wire [3:0] _GEN_334 = 4'h5 == state ? 4'h6 : _GEN_292; // @[insertSort.scala 24:19 48:19]
  wire [31:0] _GEN_335 = 4'h5 == state ? $signed(j) : $signed(_GEN_291); // @[insertSort.scala 22:16 24:19]
  wire [31:0] _GEN_336 = 4'h5 == state ? $signed(i) : $signed(_GEN_313); // @[insertSort.scala 20:16 24:19]
  wire [3:0] _GEN_337 = 4'h4 == state ? {{1'd0}, _state_T_8} : _GEN_334; // @[insertSort.scala 24:19 44:19]
  wire [31:0] _GEN_338 = 4'h4 == state ? $signed(_GEN_0) : $signed(_GEN_314); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_339 = 4'h4 == state ? $signed(_GEN_1) : $signed(_GEN_315); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_340 = 4'h4 == state ? $signed(_GEN_2) : $signed(_GEN_316); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_341 = 4'h4 == state ? $signed(_GEN_3) : $signed(_GEN_317); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_342 = 4'h4 == state ? $signed(_GEN_4) : $signed(_GEN_318); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_343 = 4'h4 == state ? $signed(_GEN_5) : $signed(_GEN_319); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_344 = 4'h4 == state ? $signed(_GEN_6) : $signed(_GEN_320); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_345 = 4'h4 == state ? $signed(_GEN_7) : $signed(_GEN_321); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_346 = 4'h4 == state ? $signed(_GEN_8) : $signed(_GEN_322); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_347 = 4'h4 == state ? $signed(_GEN_9) : $signed(_GEN_323); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_348 = 4'h4 == state ? $signed(_GEN_10) : $signed(_GEN_324); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_349 = 4'h4 == state ? $signed(_GEN_11) : $signed(_GEN_325); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_350 = 4'h4 == state ? $signed(_GEN_12) : $signed(_GEN_326); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_351 = 4'h4 == state ? $signed(_GEN_13) : $signed(_GEN_327); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_352 = 4'h4 == state ? $signed(_GEN_14) : $signed(_GEN_328); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_353 = 4'h4 == state ? $signed(_GEN_15) : $signed(_GEN_329); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_354 = 4'h4 == state ? $signed(_GEN_16) : $signed(_GEN_330); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_355 = 4'h4 == state ? $signed(_GEN_17) : $signed(_GEN_331); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_356 = 4'h4 == state ? $signed(_GEN_18) : $signed(_GEN_332); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_357 = 4'h4 == state ? $signed(_GEN_19) : $signed(_GEN_333); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_358 = 4'h4 == state ? $signed(j) : $signed(_GEN_335); // @[insertSort.scala 22:16 24:19]
  wire [31:0] _GEN_359 = 4'h4 == state ? $signed(i) : $signed(_GEN_336); // @[insertSort.scala 20:16 24:19]
  wire [31:0] _GEN_360 = 4'h3 == state ? $signed(_j_T_2) : $signed(_GEN_358); // @[insertSort.scala 24:19 40:15]
  wire [3:0] _GEN_361 = 4'h3 == state ? 4'h4 : _GEN_337; // @[insertSort.scala 24:19 41:19]
  wire [31:0] _GEN_362 = 4'h3 == state ? $signed(_GEN_0) : $signed(_GEN_338); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_363 = 4'h3 == state ? $signed(_GEN_1) : $signed(_GEN_339); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_364 = 4'h3 == state ? $signed(_GEN_2) : $signed(_GEN_340); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_365 = 4'h3 == state ? $signed(_GEN_3) : $signed(_GEN_341); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_366 = 4'h3 == state ? $signed(_GEN_4) : $signed(_GEN_342); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_367 = 4'h3 == state ? $signed(_GEN_5) : $signed(_GEN_343); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_368 = 4'h3 == state ? $signed(_GEN_6) : $signed(_GEN_344); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_369 = 4'h3 == state ? $signed(_GEN_7) : $signed(_GEN_345); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_370 = 4'h3 == state ? $signed(_GEN_8) : $signed(_GEN_346); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_371 = 4'h3 == state ? $signed(_GEN_9) : $signed(_GEN_347); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_372 = 4'h3 == state ? $signed(_GEN_10) : $signed(_GEN_348); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_373 = 4'h3 == state ? $signed(_GEN_11) : $signed(_GEN_349); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_374 = 4'h3 == state ? $signed(_GEN_12) : $signed(_GEN_350); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_375 = 4'h3 == state ? $signed(_GEN_13) : $signed(_GEN_351); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_376 = 4'h3 == state ? $signed(_GEN_14) : $signed(_GEN_352); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_377 = 4'h3 == state ? $signed(_GEN_15) : $signed(_GEN_353); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_378 = 4'h3 == state ? $signed(_GEN_16) : $signed(_GEN_354); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_379 = 4'h3 == state ? $signed(_GEN_17) : $signed(_GEN_355); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_380 = 4'h3 == state ? $signed(_GEN_18) : $signed(_GEN_356); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_381 = 4'h3 == state ? $signed(_GEN_19) : $signed(_GEN_357); // @[insertSort.scala 24:19]
  wire [31:0] _GEN_382 = 4'h3 == state ? $signed(i) : $signed(_GEN_359); // @[insertSort.scala 20:16 24:19]
  wire [3:0] _GEN_384 = 4'h2 == state ? 4'h3 : _GEN_361; // @[insertSort.scala 24:19 37:19]
  assign io_array_out_0 = array_0; // @[insertSort.scala 19:18]
  assign io_array_out_1 = array_1; // @[insertSort.scala 19:18]
  assign io_array_out_2 = array_2; // @[insertSort.scala 19:18]
  assign io_array_out_3 = array_3; // @[insertSort.scala 19:18]
  assign io_array_out_4 = array_4; // @[insertSort.scala 19:18]
  assign io_array_out_5 = array_5; // @[insertSort.scala 19:18]
  assign io_array_out_6 = array_6; // @[insertSort.scala 19:18]
  assign io_array_out_7 = array_7; // @[insertSort.scala 19:18]
  assign io_array_out_8 = array_8; // @[insertSort.scala 19:18]
  assign io_array_out_9 = array_9; // @[insertSort.scala 19:18]
  assign io_array_out_10 = array_10; // @[insertSort.scala 19:18]
  assign io_array_out_11 = array_11; // @[insertSort.scala 19:18]
  assign io_array_out_12 = array_12; // @[insertSort.scala 19:18]
  assign io_array_out_13 = array_13; // @[insertSort.scala 19:18]
  assign io_array_out_14 = array_14; // @[insertSort.scala 19:18]
  assign io_array_out_15 = array_15; // @[insertSort.scala 19:18]
  assign io_array_out_16 = array_16; // @[insertSort.scala 19:18]
  assign io_array_out_17 = array_17; // @[insertSort.scala 19:18]
  assign io_array_out_18 = array_18; // @[insertSort.scala 19:18]
  assign io_array_out_19 = array_19; // @[insertSort.scala 19:18]
  assign io_ready = state == 4'hc; // @[insertSort.scala 78:23]
  always @(posedge clock) begin
    if (reset) begin // @[insertSort.scala 13:24]
      state <= 4'hf; // @[insertSort.scala 13:24]
    end else if (4'hf == state) begin // @[insertSort.scala 24:19]
      if (io_valid) begin // @[insertSort.scala 26:25]
        state <= 4'h0;
      end
    end else if (4'h0 == state) begin // @[insertSort.scala 24:19]
      state <= 4'h1; // @[insertSort.scala 30:19]
    end else if (4'h1 == state) begin // @[insertSort.scala 24:19]
      state <= _state_T_2; // @[insertSort.scala 33:19]
    end else begin
      state <= _GEN_384;
    end
    if (4'hf == state) begin // @[insertSort.scala 24:19]
      array_0 <= _GEN_0;
    end else if (4'h0 == state) begin // @[insertSort.scala 24:19]
      array_0 <= _GEN_0;
    end else if (4'h1 == state) begin // @[insertSort.scala 24:19]
      array_0 <= _GEN_0;
    end else if (4'h2 == state) begin // @[insertSort.scala 24:19]
      array_0 <= _GEN_0;
    end else begin
      array_0 <= _GEN_362;
    end
    if (4'hf == state) begin // @[insertSort.scala 24:19]
      array_1 <= _GEN_1;
    end else if (4'h0 == state) begin // @[insertSort.scala 24:19]
      array_1 <= _GEN_1;
    end else if (4'h1 == state) begin // @[insertSort.scala 24:19]
      array_1 <= _GEN_1;
    end else if (4'h2 == state) begin // @[insertSort.scala 24:19]
      array_1 <= _GEN_1;
    end else begin
      array_1 <= _GEN_363;
    end
    if (4'hf == state) begin // @[insertSort.scala 24:19]
      array_2 <= _GEN_2;
    end else if (4'h0 == state) begin // @[insertSort.scala 24:19]
      array_2 <= _GEN_2;
    end else if (4'h1 == state) begin // @[insertSort.scala 24:19]
      array_2 <= _GEN_2;
    end else if (4'h2 == state) begin // @[insertSort.scala 24:19]
      array_2 <= _GEN_2;
    end else begin
      array_2 <= _GEN_364;
    end
    if (4'hf == state) begin // @[insertSort.scala 24:19]
      array_3 <= _GEN_3;
    end else if (4'h0 == state) begin // @[insertSort.scala 24:19]
      array_3 <= _GEN_3;
    end else if (4'h1 == state) begin // @[insertSort.scala 24:19]
      array_3 <= _GEN_3;
    end else if (4'h2 == state) begin // @[insertSort.scala 24:19]
      array_3 <= _GEN_3;
    end else begin
      array_3 <= _GEN_365;
    end
    if (4'hf == state) begin // @[insertSort.scala 24:19]
      array_4 <= _GEN_4;
    end else if (4'h0 == state) begin // @[insertSort.scala 24:19]
      array_4 <= _GEN_4;
    end else if (4'h1 == state) begin // @[insertSort.scala 24:19]
      array_4 <= _GEN_4;
    end else if (4'h2 == state) begin // @[insertSort.scala 24:19]
      array_4 <= _GEN_4;
    end else begin
      array_4 <= _GEN_366;
    end
    if (4'hf == state) begin // @[insertSort.scala 24:19]
      array_5 <= _GEN_5;
    end else if (4'h0 == state) begin // @[insertSort.scala 24:19]
      array_5 <= _GEN_5;
    end else if (4'h1 == state) begin // @[insertSort.scala 24:19]
      array_5 <= _GEN_5;
    end else if (4'h2 == state) begin // @[insertSort.scala 24:19]
      array_5 <= _GEN_5;
    end else begin
      array_5 <= _GEN_367;
    end
    if (4'hf == state) begin // @[insertSort.scala 24:19]
      array_6 <= _GEN_6;
    end else if (4'h0 == state) begin // @[insertSort.scala 24:19]
      array_6 <= _GEN_6;
    end else if (4'h1 == state) begin // @[insertSort.scala 24:19]
      array_6 <= _GEN_6;
    end else if (4'h2 == state) begin // @[insertSort.scala 24:19]
      array_6 <= _GEN_6;
    end else begin
      array_6 <= _GEN_368;
    end
    if (4'hf == state) begin // @[insertSort.scala 24:19]
      array_7 <= _GEN_7;
    end else if (4'h0 == state) begin // @[insertSort.scala 24:19]
      array_7 <= _GEN_7;
    end else if (4'h1 == state) begin // @[insertSort.scala 24:19]
      array_7 <= _GEN_7;
    end else if (4'h2 == state) begin // @[insertSort.scala 24:19]
      array_7 <= _GEN_7;
    end else begin
      array_7 <= _GEN_369;
    end
    if (4'hf == state) begin // @[insertSort.scala 24:19]
      array_8 <= _GEN_8;
    end else if (4'h0 == state) begin // @[insertSort.scala 24:19]
      array_8 <= _GEN_8;
    end else if (4'h1 == state) begin // @[insertSort.scala 24:19]
      array_8 <= _GEN_8;
    end else if (4'h2 == state) begin // @[insertSort.scala 24:19]
      array_8 <= _GEN_8;
    end else begin
      array_8 <= _GEN_370;
    end
    if (4'hf == state) begin // @[insertSort.scala 24:19]
      array_9 <= _GEN_9;
    end else if (4'h0 == state) begin // @[insertSort.scala 24:19]
      array_9 <= _GEN_9;
    end else if (4'h1 == state) begin // @[insertSort.scala 24:19]
      array_9 <= _GEN_9;
    end else if (4'h2 == state) begin // @[insertSort.scala 24:19]
      array_9 <= _GEN_9;
    end else begin
      array_9 <= _GEN_371;
    end
    if (4'hf == state) begin // @[insertSort.scala 24:19]
      array_10 <= _GEN_10;
    end else if (4'h0 == state) begin // @[insertSort.scala 24:19]
      array_10 <= _GEN_10;
    end else if (4'h1 == state) begin // @[insertSort.scala 24:19]
      array_10 <= _GEN_10;
    end else if (4'h2 == state) begin // @[insertSort.scala 24:19]
      array_10 <= _GEN_10;
    end else begin
      array_10 <= _GEN_372;
    end
    if (4'hf == state) begin // @[insertSort.scala 24:19]
      array_11 <= _GEN_11;
    end else if (4'h0 == state) begin // @[insertSort.scala 24:19]
      array_11 <= _GEN_11;
    end else if (4'h1 == state) begin // @[insertSort.scala 24:19]
      array_11 <= _GEN_11;
    end else if (4'h2 == state) begin // @[insertSort.scala 24:19]
      array_11 <= _GEN_11;
    end else begin
      array_11 <= _GEN_373;
    end
    if (4'hf == state) begin // @[insertSort.scala 24:19]
      array_12 <= _GEN_12;
    end else if (4'h0 == state) begin // @[insertSort.scala 24:19]
      array_12 <= _GEN_12;
    end else if (4'h1 == state) begin // @[insertSort.scala 24:19]
      array_12 <= _GEN_12;
    end else if (4'h2 == state) begin // @[insertSort.scala 24:19]
      array_12 <= _GEN_12;
    end else begin
      array_12 <= _GEN_374;
    end
    if (4'hf == state) begin // @[insertSort.scala 24:19]
      array_13 <= _GEN_13;
    end else if (4'h0 == state) begin // @[insertSort.scala 24:19]
      array_13 <= _GEN_13;
    end else if (4'h1 == state) begin // @[insertSort.scala 24:19]
      array_13 <= _GEN_13;
    end else if (4'h2 == state) begin // @[insertSort.scala 24:19]
      array_13 <= _GEN_13;
    end else begin
      array_13 <= _GEN_375;
    end
    if (4'hf == state) begin // @[insertSort.scala 24:19]
      array_14 <= _GEN_14;
    end else if (4'h0 == state) begin // @[insertSort.scala 24:19]
      array_14 <= _GEN_14;
    end else if (4'h1 == state) begin // @[insertSort.scala 24:19]
      array_14 <= _GEN_14;
    end else if (4'h2 == state) begin // @[insertSort.scala 24:19]
      array_14 <= _GEN_14;
    end else begin
      array_14 <= _GEN_376;
    end
    if (4'hf == state) begin // @[insertSort.scala 24:19]
      array_15 <= _GEN_15;
    end else if (4'h0 == state) begin // @[insertSort.scala 24:19]
      array_15 <= _GEN_15;
    end else if (4'h1 == state) begin // @[insertSort.scala 24:19]
      array_15 <= _GEN_15;
    end else if (4'h2 == state) begin // @[insertSort.scala 24:19]
      array_15 <= _GEN_15;
    end else begin
      array_15 <= _GEN_377;
    end
    if (4'hf == state) begin // @[insertSort.scala 24:19]
      array_16 <= _GEN_16;
    end else if (4'h0 == state) begin // @[insertSort.scala 24:19]
      array_16 <= _GEN_16;
    end else if (4'h1 == state) begin // @[insertSort.scala 24:19]
      array_16 <= _GEN_16;
    end else if (4'h2 == state) begin // @[insertSort.scala 24:19]
      array_16 <= _GEN_16;
    end else begin
      array_16 <= _GEN_378;
    end
    if (4'hf == state) begin // @[insertSort.scala 24:19]
      array_17 <= _GEN_17;
    end else if (4'h0 == state) begin // @[insertSort.scala 24:19]
      array_17 <= _GEN_17;
    end else if (4'h1 == state) begin // @[insertSort.scala 24:19]
      array_17 <= _GEN_17;
    end else if (4'h2 == state) begin // @[insertSort.scala 24:19]
      array_17 <= _GEN_17;
    end else begin
      array_17 <= _GEN_379;
    end
    if (4'hf == state) begin // @[insertSort.scala 24:19]
      array_18 <= _GEN_18;
    end else if (4'h0 == state) begin // @[insertSort.scala 24:19]
      array_18 <= _GEN_18;
    end else if (4'h1 == state) begin // @[insertSort.scala 24:19]
      array_18 <= _GEN_18;
    end else if (4'h2 == state) begin // @[insertSort.scala 24:19]
      array_18 <= _GEN_18;
    end else begin
      array_18 <= _GEN_380;
    end
    if (4'hf == state) begin // @[insertSort.scala 24:19]
      array_19 <= _GEN_19;
    end else if (4'h0 == state) begin // @[insertSort.scala 24:19]
      array_19 <= _GEN_19;
    end else if (4'h1 == state) begin // @[insertSort.scala 24:19]
      array_19 <= _GEN_19;
    end else if (4'h2 == state) begin // @[insertSort.scala 24:19]
      array_19 <= _GEN_19;
    end else begin
      array_19 <= _GEN_381;
    end
    REG <= ~io_valid; // @[insertSort.scala 16:18]
    if (!(4'hf == state)) begin // @[insertSort.scala 24:19]
      if (4'h0 == state) begin // @[insertSort.scala 24:19]
        i <= 32'sh1; // @[insertSort.scala 29:15]
      end else if (!(4'h1 == state)) begin // @[insertSort.scala 24:19]
        if (!(4'h2 == state)) begin // @[insertSort.scala 24:19]
          i <= _GEN_382;
        end
      end
    end
    if (!(4'hf == state)) begin // @[insertSort.scala 24:19]
      if (!(4'h0 == state)) begin // @[insertSort.scala 24:19]
        if (!(4'h1 == state)) begin // @[insertSort.scala 24:19]
          if (4'h2 == state) begin // @[insertSort.scala 24:19]
            key <= _GEN_39; // @[insertSort.scala 36:17]
          end
        end
      end
    end
    if (!(4'hf == state)) begin // @[insertSort.scala 24:19]
      if (!(4'h0 == state)) begin // @[insertSort.scala 24:19]
        if (!(4'h1 == state)) begin // @[insertSort.scala 24:19]
          if (!(4'h2 == state)) begin // @[insertSort.scala 24:19]
            j <= _GEN_360;
          end
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  array_0 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  array_1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  array_2 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  array_3 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  array_4 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  array_5 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  array_6 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  array_7 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  array_8 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  array_9 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  array_10 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  array_11 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  array_12 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  array_13 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  array_14 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  array_15 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  array_16 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  array_17 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  array_18 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  array_19 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  REG = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  i = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  key = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  j = _RAND_24[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
